* Example 01 SPICE subckt definition

.subckt example_01 input[1] input[0] output[0] input[2] control
* Circuit internals omitted
.ends
