* circuit.Package sramgen_sramgen_sram_128x64m2w64_replica_v1
* Written by SpiceNetlister
* 

.SUBCKT hierarchical_decoder_nand_2 
+ gnd vdd a b c y 

xn1 
+ x1 a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ x2 b x1 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn3 
+ y c x2 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp3 
+ y c vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder_inv_3 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder_nand_53 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder 
+ vdd gnd addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] addr_b[5] addr_b[4] addr_b[3] addr_b[2] addr_b[1] addr_b[0] decode[63] decode[62] decode[61] decode[60] decode[59] decode[58] decode[57] decode[56] decode[55] decode[54] decode[53] decode[52] decode[51] decode[50] decode[49] decode[48] decode[47] decode[46] decode[45] decode[44] decode[43] decode[42] decode[41] decode[40] decode[39] decode[38] decode[37] decode[36] decode[35] decode[34] decode[33] decode[32] decode[31] decode[30] decode[29] decode[28] decode[27] decode[26] decode[25] decode[24] decode[23] decode[22] decode[21] decode[20] decode[19] decode[18] decode[17] decode[16] decode[15] decode[14] decode[13] decode[12] decode[11] decode[10] decode[9] decode[8] decode[7] decode[6] decode[5] decode[4] decode[3] decode[2] decode[1] decode[0] decode_b[63] decode_b[62] decode_b[61] decode_b[60] decode_b[59] decode_b[58] decode_b[57] decode_b[56] decode_b[55] decode_b[54] decode_b[53] decode_b[52] decode_b[51] decode_b[50] decode_b[49] decode_b[48] decode_b[47] decode_b[46] decode_b[45] decode_b[44] decode_b[43] decode_b[42] decode_b[41] decode_b[40] decode_b[39] decode_b[38] decode_b[37] decode_b[36] decode_b[35] decode_b[34] decode_b[33] decode_b[32] decode_b[31] decode_b[30] decode_b[29] decode_b[28] decode_b[27] decode_b[26] decode_b[25] decode_b[24] decode_b[23] decode_b[22] decode_b[21] decode_b[20] decode_b[19] decode_b[18] decode_b[17] decode_b[16] decode_b[15] decode_b[14] decode_b[13] decode_b[12] decode_b[11] decode_b[10] decode_b[9] decode_b[8] decode_b[7] decode_b[6] decode_b[5] decode_b[4] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_5 
+ gnd vdd addr_b[5] addr_b[4] addr_b[3] net_4 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_6 
+ gnd vdd net_4 predecode_1[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_8 
+ gnd vdd addr_b[5] addr_b[4] addr[3] net_7 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_9 
+ gnd vdd net_7 predecode_1[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_11 
+ gnd vdd addr_b[5] addr[4] addr_b[3] net_10 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_12 
+ gnd vdd net_10 predecode_1[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_14 
+ gnd vdd addr_b[5] addr[4] addr[3] net_13 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_15 
+ gnd vdd net_13 predecode_1[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_17 
+ gnd vdd addr[5] addr_b[4] addr_b[3] net_16 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_18 
+ gnd vdd net_16 predecode_1[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_20 
+ gnd vdd addr[5] addr_b[4] addr[3] net_19 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_21 
+ gnd vdd net_19 predecode_1[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_23 
+ gnd vdd addr[5] addr[4] addr_b[3] net_22 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_24 
+ gnd vdd net_22 predecode_1[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_26 
+ gnd vdd addr[5] addr[4] addr[3] net_25 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_27 
+ gnd vdd net_25 predecode_1[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_30 
+ gnd vdd addr_b[2] addr_b[1] addr_b[0] net_29 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_31 
+ gnd vdd net_29 predecode_28[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_33 
+ gnd vdd addr_b[2] addr_b[1] addr[0] net_32 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_34 
+ gnd vdd net_32 predecode_28[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_36 
+ gnd vdd addr_b[2] addr[1] addr_b[0] net_35 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_37 
+ gnd vdd net_35 predecode_28[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_39 
+ gnd vdd addr_b[2] addr[1] addr[0] net_38 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_40 
+ gnd vdd net_38 predecode_28[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_42 
+ gnd vdd addr[2] addr_b[1] addr_b[0] net_41 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_43 
+ gnd vdd net_41 predecode_28[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_45 
+ gnd vdd addr[2] addr_b[1] addr[0] net_44 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_46 
+ gnd vdd net_44 predecode_28[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_48 
+ gnd vdd addr[2] addr[1] addr_b[0] net_47 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_49 
+ gnd vdd net_47 predecode_28[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_51 
+ gnd vdd addr[2] addr[1] addr[0] net_50 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_52 
+ gnd vdd net_50 predecode_28[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_54 
+ gnd vdd predecode_1[0] predecode_28[0] decode_b[0] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_55 
+ gnd vdd decode_b[0] decode[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_56 
+ gnd vdd predecode_1[0] predecode_28[1] decode_b[1] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_57 
+ gnd vdd decode_b[1] decode[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_58 
+ gnd vdd predecode_1[0] predecode_28[2] decode_b[2] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_59 
+ gnd vdd decode_b[2] decode[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_60 
+ gnd vdd predecode_1[0] predecode_28[3] decode_b[3] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_61 
+ gnd vdd decode_b[3] decode[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_62 
+ gnd vdd predecode_1[0] predecode_28[4] decode_b[4] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_63 
+ gnd vdd decode_b[4] decode[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_64 
+ gnd vdd predecode_1[0] predecode_28[5] decode_b[5] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_65 
+ gnd vdd decode_b[5] decode[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_66 
+ gnd vdd predecode_1[0] predecode_28[6] decode_b[6] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_67 
+ gnd vdd decode_b[6] decode[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_68 
+ gnd vdd predecode_1[0] predecode_28[7] decode_b[7] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_69 
+ gnd vdd decode_b[7] decode[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_70 
+ gnd vdd predecode_1[1] predecode_28[0] decode_b[8] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_71 
+ gnd vdd decode_b[8] decode[8] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_72 
+ gnd vdd predecode_1[1] predecode_28[1] decode_b[9] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_73 
+ gnd vdd decode_b[9] decode[9] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_74 
+ gnd vdd predecode_1[1] predecode_28[2] decode_b[10] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_75 
+ gnd vdd decode_b[10] decode[10] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_76 
+ gnd vdd predecode_1[1] predecode_28[3] decode_b[11] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_77 
+ gnd vdd decode_b[11] decode[11] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_78 
+ gnd vdd predecode_1[1] predecode_28[4] decode_b[12] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_79 
+ gnd vdd decode_b[12] decode[12] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_80 
+ gnd vdd predecode_1[1] predecode_28[5] decode_b[13] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_81 
+ gnd vdd decode_b[13] decode[13] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_82 
+ gnd vdd predecode_1[1] predecode_28[6] decode_b[14] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_83 
+ gnd vdd decode_b[14] decode[14] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_84 
+ gnd vdd predecode_1[1] predecode_28[7] decode_b[15] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_85 
+ gnd vdd decode_b[15] decode[15] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_86 
+ gnd vdd predecode_1[2] predecode_28[0] decode_b[16] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_87 
+ gnd vdd decode_b[16] decode[16] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_88 
+ gnd vdd predecode_1[2] predecode_28[1] decode_b[17] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_89 
+ gnd vdd decode_b[17] decode[17] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_90 
+ gnd vdd predecode_1[2] predecode_28[2] decode_b[18] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_91 
+ gnd vdd decode_b[18] decode[18] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_92 
+ gnd vdd predecode_1[2] predecode_28[3] decode_b[19] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_93 
+ gnd vdd decode_b[19] decode[19] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_94 
+ gnd vdd predecode_1[2] predecode_28[4] decode_b[20] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_95 
+ gnd vdd decode_b[20] decode[20] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_96 
+ gnd vdd predecode_1[2] predecode_28[5] decode_b[21] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_97 
+ gnd vdd decode_b[21] decode[21] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_98 
+ gnd vdd predecode_1[2] predecode_28[6] decode_b[22] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_99 
+ gnd vdd decode_b[22] decode[22] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_100 
+ gnd vdd predecode_1[2] predecode_28[7] decode_b[23] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_101 
+ gnd vdd decode_b[23] decode[23] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_102 
+ gnd vdd predecode_1[3] predecode_28[0] decode_b[24] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_103 
+ gnd vdd decode_b[24] decode[24] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_104 
+ gnd vdd predecode_1[3] predecode_28[1] decode_b[25] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_105 
+ gnd vdd decode_b[25] decode[25] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_106 
+ gnd vdd predecode_1[3] predecode_28[2] decode_b[26] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_107 
+ gnd vdd decode_b[26] decode[26] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_108 
+ gnd vdd predecode_1[3] predecode_28[3] decode_b[27] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_109 
+ gnd vdd decode_b[27] decode[27] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_110 
+ gnd vdd predecode_1[3] predecode_28[4] decode_b[28] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_111 
+ gnd vdd decode_b[28] decode[28] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_112 
+ gnd vdd predecode_1[3] predecode_28[5] decode_b[29] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_113 
+ gnd vdd decode_b[29] decode[29] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_114 
+ gnd vdd predecode_1[3] predecode_28[6] decode_b[30] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_115 
+ gnd vdd decode_b[30] decode[30] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_116 
+ gnd vdd predecode_1[3] predecode_28[7] decode_b[31] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_117 
+ gnd vdd decode_b[31] decode[31] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_118 
+ gnd vdd predecode_1[4] predecode_28[0] decode_b[32] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_119 
+ gnd vdd decode_b[32] decode[32] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_120 
+ gnd vdd predecode_1[4] predecode_28[1] decode_b[33] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_121 
+ gnd vdd decode_b[33] decode[33] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_122 
+ gnd vdd predecode_1[4] predecode_28[2] decode_b[34] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_123 
+ gnd vdd decode_b[34] decode[34] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_124 
+ gnd vdd predecode_1[4] predecode_28[3] decode_b[35] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_125 
+ gnd vdd decode_b[35] decode[35] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_126 
+ gnd vdd predecode_1[4] predecode_28[4] decode_b[36] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_127 
+ gnd vdd decode_b[36] decode[36] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_128 
+ gnd vdd predecode_1[4] predecode_28[5] decode_b[37] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_129 
+ gnd vdd decode_b[37] decode[37] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_130 
+ gnd vdd predecode_1[4] predecode_28[6] decode_b[38] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_131 
+ gnd vdd decode_b[38] decode[38] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_132 
+ gnd vdd predecode_1[4] predecode_28[7] decode_b[39] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_133 
+ gnd vdd decode_b[39] decode[39] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_134 
+ gnd vdd predecode_1[5] predecode_28[0] decode_b[40] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_135 
+ gnd vdd decode_b[40] decode[40] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_136 
+ gnd vdd predecode_1[5] predecode_28[1] decode_b[41] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_137 
+ gnd vdd decode_b[41] decode[41] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_138 
+ gnd vdd predecode_1[5] predecode_28[2] decode_b[42] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_139 
+ gnd vdd decode_b[42] decode[42] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_140 
+ gnd vdd predecode_1[5] predecode_28[3] decode_b[43] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_141 
+ gnd vdd decode_b[43] decode[43] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_142 
+ gnd vdd predecode_1[5] predecode_28[4] decode_b[44] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_143 
+ gnd vdd decode_b[44] decode[44] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_144 
+ gnd vdd predecode_1[5] predecode_28[5] decode_b[45] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_145 
+ gnd vdd decode_b[45] decode[45] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_146 
+ gnd vdd predecode_1[5] predecode_28[6] decode_b[46] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_147 
+ gnd vdd decode_b[46] decode[46] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_148 
+ gnd vdd predecode_1[5] predecode_28[7] decode_b[47] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_149 
+ gnd vdd decode_b[47] decode[47] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_150 
+ gnd vdd predecode_1[6] predecode_28[0] decode_b[48] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_151 
+ gnd vdd decode_b[48] decode[48] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_152 
+ gnd vdd predecode_1[6] predecode_28[1] decode_b[49] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_153 
+ gnd vdd decode_b[49] decode[49] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_154 
+ gnd vdd predecode_1[6] predecode_28[2] decode_b[50] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_155 
+ gnd vdd decode_b[50] decode[50] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_156 
+ gnd vdd predecode_1[6] predecode_28[3] decode_b[51] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_157 
+ gnd vdd decode_b[51] decode[51] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_158 
+ gnd vdd predecode_1[6] predecode_28[4] decode_b[52] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_159 
+ gnd vdd decode_b[52] decode[52] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_160 
+ gnd vdd predecode_1[6] predecode_28[5] decode_b[53] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_161 
+ gnd vdd decode_b[53] decode[53] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_162 
+ gnd vdd predecode_1[6] predecode_28[6] decode_b[54] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_163 
+ gnd vdd decode_b[54] decode[54] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_164 
+ gnd vdd predecode_1[6] predecode_28[7] decode_b[55] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_165 
+ gnd vdd decode_b[55] decode[55] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_166 
+ gnd vdd predecode_1[7] predecode_28[0] decode_b[56] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_167 
+ gnd vdd decode_b[56] decode[56] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_168 
+ gnd vdd predecode_1[7] predecode_28[1] decode_b[57] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_169 
+ gnd vdd decode_b[57] decode[57] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_170 
+ gnd vdd predecode_1[7] predecode_28[2] decode_b[58] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_171 
+ gnd vdd decode_b[58] decode[58] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_172 
+ gnd vdd predecode_1[7] predecode_28[3] decode_b[59] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_173 
+ gnd vdd decode_b[59] decode[59] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_174 
+ gnd vdd predecode_1[7] predecode_28[4] decode_b[60] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_175 
+ gnd vdd decode_b[60] decode[60] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_176 
+ gnd vdd predecode_1[7] predecode_28[5] decode_b[61] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_177 
+ gnd vdd decode_b[61] decode[61] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_178 
+ gnd vdd predecode_1[7] predecode_28[6] decode_b[62] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_179 
+ gnd vdd decode_b[62] decode[62] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_180 
+ gnd vdd predecode_1[7] predecode_28[7] decode_b[63] 
+ hierarchical_decoder_nand_53 
* No parameters

xinv_181 
+ gnd vdd decode_b[63] decode[63] 
+ hierarchical_decoder_inv_3 
* No parameters

.ENDS

.SUBCKT wordline_driver_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ wordline_driver_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ wordline_driver_and2_inv 
* No parameters

.ENDS

.SUBCKT wordline_driver 
+ vdd vss din wl_en wl 

xand2 
+ din wl_en wl vdd vss 
+ wordline_driver_and2 
* No parameters

.ENDS

.SUBCKT wordline_driver_array 
+ vdd vss din[63] din[62] din[61] din[60] din[59] din[58] din[57] din[56] din[55] din[54] din[53] din[52] din[51] din[50] din[49] din[48] din[47] din[46] din[45] din[44] din[43] din[42] din[41] din[40] din[39] din[38] din[37] din[36] din[35] din[34] din[33] din[32] din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] wl_en wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] 

xwl_driver_0 
+ vdd vss din[0] wl_en wl[0] 
+ wordline_driver 
* No parameters

xwl_driver_1 
+ vdd vss din[1] wl_en wl[1] 
+ wordline_driver 
* No parameters

xwl_driver_2 
+ vdd vss din[2] wl_en wl[2] 
+ wordline_driver 
* No parameters

xwl_driver_3 
+ vdd vss din[3] wl_en wl[3] 
+ wordline_driver 
* No parameters

xwl_driver_4 
+ vdd vss din[4] wl_en wl[4] 
+ wordline_driver 
* No parameters

xwl_driver_5 
+ vdd vss din[5] wl_en wl[5] 
+ wordline_driver 
* No parameters

xwl_driver_6 
+ vdd vss din[6] wl_en wl[6] 
+ wordline_driver 
* No parameters

xwl_driver_7 
+ vdd vss din[7] wl_en wl[7] 
+ wordline_driver 
* No parameters

xwl_driver_8 
+ vdd vss din[8] wl_en wl[8] 
+ wordline_driver 
* No parameters

xwl_driver_9 
+ vdd vss din[9] wl_en wl[9] 
+ wordline_driver 
* No parameters

xwl_driver_10 
+ vdd vss din[10] wl_en wl[10] 
+ wordline_driver 
* No parameters

xwl_driver_11 
+ vdd vss din[11] wl_en wl[11] 
+ wordline_driver 
* No parameters

xwl_driver_12 
+ vdd vss din[12] wl_en wl[12] 
+ wordline_driver 
* No parameters

xwl_driver_13 
+ vdd vss din[13] wl_en wl[13] 
+ wordline_driver 
* No parameters

xwl_driver_14 
+ vdd vss din[14] wl_en wl[14] 
+ wordline_driver 
* No parameters

xwl_driver_15 
+ vdd vss din[15] wl_en wl[15] 
+ wordline_driver 
* No parameters

xwl_driver_16 
+ vdd vss din[16] wl_en wl[16] 
+ wordline_driver 
* No parameters

xwl_driver_17 
+ vdd vss din[17] wl_en wl[17] 
+ wordline_driver 
* No parameters

xwl_driver_18 
+ vdd vss din[18] wl_en wl[18] 
+ wordline_driver 
* No parameters

xwl_driver_19 
+ vdd vss din[19] wl_en wl[19] 
+ wordline_driver 
* No parameters

xwl_driver_20 
+ vdd vss din[20] wl_en wl[20] 
+ wordline_driver 
* No parameters

xwl_driver_21 
+ vdd vss din[21] wl_en wl[21] 
+ wordline_driver 
* No parameters

xwl_driver_22 
+ vdd vss din[22] wl_en wl[22] 
+ wordline_driver 
* No parameters

xwl_driver_23 
+ vdd vss din[23] wl_en wl[23] 
+ wordline_driver 
* No parameters

xwl_driver_24 
+ vdd vss din[24] wl_en wl[24] 
+ wordline_driver 
* No parameters

xwl_driver_25 
+ vdd vss din[25] wl_en wl[25] 
+ wordline_driver 
* No parameters

xwl_driver_26 
+ vdd vss din[26] wl_en wl[26] 
+ wordline_driver 
* No parameters

xwl_driver_27 
+ vdd vss din[27] wl_en wl[27] 
+ wordline_driver 
* No parameters

xwl_driver_28 
+ vdd vss din[28] wl_en wl[28] 
+ wordline_driver 
* No parameters

xwl_driver_29 
+ vdd vss din[29] wl_en wl[29] 
+ wordline_driver 
* No parameters

xwl_driver_30 
+ vdd vss din[30] wl_en wl[30] 
+ wordline_driver 
* No parameters

xwl_driver_31 
+ vdd vss din[31] wl_en wl[31] 
+ wordline_driver 
* No parameters

xwl_driver_32 
+ vdd vss din[32] wl_en wl[32] 
+ wordline_driver 
* No parameters

xwl_driver_33 
+ vdd vss din[33] wl_en wl[33] 
+ wordline_driver 
* No parameters

xwl_driver_34 
+ vdd vss din[34] wl_en wl[34] 
+ wordline_driver 
* No parameters

xwl_driver_35 
+ vdd vss din[35] wl_en wl[35] 
+ wordline_driver 
* No parameters

xwl_driver_36 
+ vdd vss din[36] wl_en wl[36] 
+ wordline_driver 
* No parameters

xwl_driver_37 
+ vdd vss din[37] wl_en wl[37] 
+ wordline_driver 
* No parameters

xwl_driver_38 
+ vdd vss din[38] wl_en wl[38] 
+ wordline_driver 
* No parameters

xwl_driver_39 
+ vdd vss din[39] wl_en wl[39] 
+ wordline_driver 
* No parameters

xwl_driver_40 
+ vdd vss din[40] wl_en wl[40] 
+ wordline_driver 
* No parameters

xwl_driver_41 
+ vdd vss din[41] wl_en wl[41] 
+ wordline_driver 
* No parameters

xwl_driver_42 
+ vdd vss din[42] wl_en wl[42] 
+ wordline_driver 
* No parameters

xwl_driver_43 
+ vdd vss din[43] wl_en wl[43] 
+ wordline_driver 
* No parameters

xwl_driver_44 
+ vdd vss din[44] wl_en wl[44] 
+ wordline_driver 
* No parameters

xwl_driver_45 
+ vdd vss din[45] wl_en wl[45] 
+ wordline_driver 
* No parameters

xwl_driver_46 
+ vdd vss din[46] wl_en wl[46] 
+ wordline_driver 
* No parameters

xwl_driver_47 
+ vdd vss din[47] wl_en wl[47] 
+ wordline_driver 
* No parameters

xwl_driver_48 
+ vdd vss din[48] wl_en wl[48] 
+ wordline_driver 
* No parameters

xwl_driver_49 
+ vdd vss din[49] wl_en wl[49] 
+ wordline_driver 
* No parameters

xwl_driver_50 
+ vdd vss din[50] wl_en wl[50] 
+ wordline_driver 
* No parameters

xwl_driver_51 
+ vdd vss din[51] wl_en wl[51] 
+ wordline_driver 
* No parameters

xwl_driver_52 
+ vdd vss din[52] wl_en wl[52] 
+ wordline_driver 
* No parameters

xwl_driver_53 
+ vdd vss din[53] wl_en wl[53] 
+ wordline_driver 
* No parameters

xwl_driver_54 
+ vdd vss din[54] wl_en wl[54] 
+ wordline_driver 
* No parameters

xwl_driver_55 
+ vdd vss din[55] wl_en wl[55] 
+ wordline_driver 
* No parameters

xwl_driver_56 
+ vdd vss din[56] wl_en wl[56] 
+ wordline_driver 
* No parameters

xwl_driver_57 
+ vdd vss din[57] wl_en wl[57] 
+ wordline_driver 
* No parameters

xwl_driver_58 
+ vdd vss din[58] wl_en wl[58] 
+ wordline_driver 
* No parameters

xwl_driver_59 
+ vdd vss din[59] wl_en wl[59] 
+ wordline_driver 
* No parameters

xwl_driver_60 
+ vdd vss din[60] wl_en wl[60] 
+ wordline_driver 
* No parameters

xwl_driver_61 
+ vdd vss din[61] wl_en wl[61] 
+ wordline_driver 
* No parameters

xwl_driver_62 
+ vdd vss din[62] wl_en wl[62] 
+ wordline_driver 
* No parameters

xwl_driver_63 
+ vdd vss din[63] wl_en wl[63] 
+ wordline_driver 
* No parameters

.ENDS

.SUBCKT bitcell_array 
+ vdd vss bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] vnb vpb rbl rbr 

xbitcell_0_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_130 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_131 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_130 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_131 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_0 
+ vdd vdd vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_1 
+ rbl rbr vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_2 
+ bl[0] br[0] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_3 
+ bl[1] br[1] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_4 
+ bl[2] br[2] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_5 
+ bl[3] br[3] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_6 
+ bl[4] br[4] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_7 
+ bl[5] br[5] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_8 
+ bl[6] br[6] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_9 
+ bl[7] br[7] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_10 
+ bl[8] br[8] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_11 
+ bl[9] br[9] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_12 
+ bl[10] br[10] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_13 
+ bl[11] br[11] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_14 
+ bl[12] br[12] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_15 
+ bl[13] br[13] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_16 
+ bl[14] br[14] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_17 
+ bl[15] br[15] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_18 
+ bl[16] br[16] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_19 
+ bl[17] br[17] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_20 
+ bl[18] br[18] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_21 
+ bl[19] br[19] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_22 
+ bl[20] br[20] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_23 
+ bl[21] br[21] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_24 
+ bl[22] br[22] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_25 
+ bl[23] br[23] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_26 
+ bl[24] br[24] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_27 
+ bl[25] br[25] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_28 
+ bl[26] br[26] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_29 
+ bl[27] br[27] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_30 
+ bl[28] br[28] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_31 
+ bl[29] br[29] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_32 
+ bl[30] br[30] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_33 
+ bl[31] br[31] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_34 
+ bl[32] br[32] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_35 
+ bl[33] br[33] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_36 
+ bl[34] br[34] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_37 
+ bl[35] br[35] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_38 
+ bl[36] br[36] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_39 
+ bl[37] br[37] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_40 
+ bl[38] br[38] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_41 
+ bl[39] br[39] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_42 
+ bl[40] br[40] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_43 
+ bl[41] br[41] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_44 
+ bl[42] br[42] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_45 
+ bl[43] br[43] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_46 
+ bl[44] br[44] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_47 
+ bl[45] br[45] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_48 
+ bl[46] br[46] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_49 
+ bl[47] br[47] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_50 
+ bl[48] br[48] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_51 
+ bl[49] br[49] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_52 
+ bl[50] br[50] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_53 
+ bl[51] br[51] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_54 
+ bl[52] br[52] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_55 
+ bl[53] br[53] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_56 
+ bl[54] br[54] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_57 
+ bl[55] br[55] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_58 
+ bl[56] br[56] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_59 
+ bl[57] br[57] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_60 
+ bl[58] br[58] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_61 
+ bl[59] br[59] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_62 
+ bl[60] br[60] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_63 
+ bl[61] br[61] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_64 
+ bl[62] br[62] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_65 
+ bl[63] br[63] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_66 
+ bl[64] br[64] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_67 
+ bl[65] br[65] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_68 
+ bl[66] br[66] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_69 
+ bl[67] br[67] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_70 
+ bl[68] br[68] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_71 
+ bl[69] br[69] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_72 
+ bl[70] br[70] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_73 
+ bl[71] br[71] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_74 
+ bl[72] br[72] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_75 
+ bl[73] br[73] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_76 
+ bl[74] br[74] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_77 
+ bl[75] br[75] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_78 
+ bl[76] br[76] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_79 
+ bl[77] br[77] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_80 
+ bl[78] br[78] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_81 
+ bl[79] br[79] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_82 
+ bl[80] br[80] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_83 
+ bl[81] br[81] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_84 
+ bl[82] br[82] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_85 
+ bl[83] br[83] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_86 
+ bl[84] br[84] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_87 
+ bl[85] br[85] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_88 
+ bl[86] br[86] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_89 
+ bl[87] br[87] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_90 
+ bl[88] br[88] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_91 
+ bl[89] br[89] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_92 
+ bl[90] br[90] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_93 
+ bl[91] br[91] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_94 
+ bl[92] br[92] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_95 
+ bl[93] br[93] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_96 
+ bl[94] br[94] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_97 
+ bl[95] br[95] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_98 
+ bl[96] br[96] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_99 
+ bl[97] br[97] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_100 
+ bl[98] br[98] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_101 
+ bl[99] br[99] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_102 
+ bl[100] br[100] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_103 
+ bl[101] br[101] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_104 
+ bl[102] br[102] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_105 
+ bl[103] br[103] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_106 
+ bl[104] br[104] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_107 
+ bl[105] br[105] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_108 
+ bl[106] br[106] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_109 
+ bl[107] br[107] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_110 
+ bl[108] br[108] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_111 
+ bl[109] br[109] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_112 
+ bl[110] br[110] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_113 
+ bl[111] br[111] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_114 
+ bl[112] br[112] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_115 
+ bl[113] br[113] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_116 
+ bl[114] br[114] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_117 
+ bl[115] br[115] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_118 
+ bl[116] br[116] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_119 
+ bl[117] br[117] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_120 
+ bl[118] br[118] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_121 
+ bl[119] br[119] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_122 
+ bl[120] br[120] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_123 
+ bl[121] br[121] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_124 
+ bl[122] br[122] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_125 
+ bl[123] br[123] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_126 
+ bl[124] br[124] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_127 
+ bl[125] br[125] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_128 
+ bl[126] br[126] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_129 
+ bl[127] br[127] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_130 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_131 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_0 
+ vdd vdd vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_1 
+ rbl rbr vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_2 
+ bl[0] br[0] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_3 
+ bl[1] br[1] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_4 
+ bl[2] br[2] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_5 
+ bl[3] br[3] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_6 
+ bl[4] br[4] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_7 
+ bl[5] br[5] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_8 
+ bl[6] br[6] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_9 
+ bl[7] br[7] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_10 
+ bl[8] br[8] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_11 
+ bl[9] br[9] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_12 
+ bl[10] br[10] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_13 
+ bl[11] br[11] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_14 
+ bl[12] br[12] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_15 
+ bl[13] br[13] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_16 
+ bl[14] br[14] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_17 
+ bl[15] br[15] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_18 
+ bl[16] br[16] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_19 
+ bl[17] br[17] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_20 
+ bl[18] br[18] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_21 
+ bl[19] br[19] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_22 
+ bl[20] br[20] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_23 
+ bl[21] br[21] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_24 
+ bl[22] br[22] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_25 
+ bl[23] br[23] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_26 
+ bl[24] br[24] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_27 
+ bl[25] br[25] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_28 
+ bl[26] br[26] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_29 
+ bl[27] br[27] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_30 
+ bl[28] br[28] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_31 
+ bl[29] br[29] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_32 
+ bl[30] br[30] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_33 
+ bl[31] br[31] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_34 
+ bl[32] br[32] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_35 
+ bl[33] br[33] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_36 
+ bl[34] br[34] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_37 
+ bl[35] br[35] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_38 
+ bl[36] br[36] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_39 
+ bl[37] br[37] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_40 
+ bl[38] br[38] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_41 
+ bl[39] br[39] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_42 
+ bl[40] br[40] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_43 
+ bl[41] br[41] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_44 
+ bl[42] br[42] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_45 
+ bl[43] br[43] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_46 
+ bl[44] br[44] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_47 
+ bl[45] br[45] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_48 
+ bl[46] br[46] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_49 
+ bl[47] br[47] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_50 
+ bl[48] br[48] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_51 
+ bl[49] br[49] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_52 
+ bl[50] br[50] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_53 
+ bl[51] br[51] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_54 
+ bl[52] br[52] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_55 
+ bl[53] br[53] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_56 
+ bl[54] br[54] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_57 
+ bl[55] br[55] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_58 
+ bl[56] br[56] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_59 
+ bl[57] br[57] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_60 
+ bl[58] br[58] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_61 
+ bl[59] br[59] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_62 
+ bl[60] br[60] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_63 
+ bl[61] br[61] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_64 
+ bl[62] br[62] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_65 
+ bl[63] br[63] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_66 
+ bl[64] br[64] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_67 
+ bl[65] br[65] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_68 
+ bl[66] br[66] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_69 
+ bl[67] br[67] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_70 
+ bl[68] br[68] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_71 
+ bl[69] br[69] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_72 
+ bl[70] br[70] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_73 
+ bl[71] br[71] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_74 
+ bl[72] br[72] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_75 
+ bl[73] br[73] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_76 
+ bl[74] br[74] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_77 
+ bl[75] br[75] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_78 
+ bl[76] br[76] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_79 
+ bl[77] br[77] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_80 
+ bl[78] br[78] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_81 
+ bl[79] br[79] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_82 
+ bl[80] br[80] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_83 
+ bl[81] br[81] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_84 
+ bl[82] br[82] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_85 
+ bl[83] br[83] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_86 
+ bl[84] br[84] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_87 
+ bl[85] br[85] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_88 
+ bl[86] br[86] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_89 
+ bl[87] br[87] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_90 
+ bl[88] br[88] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_91 
+ bl[89] br[89] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_92 
+ bl[90] br[90] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_93 
+ bl[91] br[91] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_94 
+ bl[92] br[92] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_95 
+ bl[93] br[93] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_96 
+ bl[94] br[94] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_97 
+ bl[95] br[95] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_98 
+ bl[96] br[96] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_99 
+ bl[97] br[97] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_100 
+ bl[98] br[98] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_101 
+ bl[99] br[99] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_102 
+ bl[100] br[100] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_103 
+ bl[101] br[101] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_104 
+ bl[102] br[102] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_105 
+ bl[103] br[103] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_106 
+ bl[104] br[104] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_107 
+ bl[105] br[105] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_108 
+ bl[106] br[106] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_109 
+ bl[107] br[107] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_110 
+ bl[108] br[108] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_111 
+ bl[109] br[109] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_112 
+ bl[110] br[110] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_113 
+ bl[111] br[111] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_114 
+ bl[112] br[112] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_115 
+ bl[113] br[113] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_116 
+ bl[114] br[114] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_117 
+ bl[115] br[115] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_118 
+ bl[116] br[116] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_119 
+ bl[117] br[117] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_120 
+ bl[118] br[118] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_121 
+ bl[119] br[119] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_122 
+ bl[120] br[120] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_123 
+ bl[121] br[121] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_124 
+ bl[122] br[122] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_125 
+ bl[123] br[123] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_126 
+ bl[124] br[124] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_127 
+ bl[125] br[125] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_128 
+ bl[126] br[126] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_129 
+ bl[127] br[127] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_130 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_131 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_0 
+ vdd vdd vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_1 
+ rbl rbr vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_2 
+ bl[0] br[0] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_3 
+ bl[1] br[1] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_4 
+ bl[2] br[2] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_5 
+ bl[3] br[3] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_6 
+ bl[4] br[4] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_7 
+ bl[5] br[5] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_8 
+ bl[6] br[6] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_9 
+ bl[7] br[7] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_10 
+ bl[8] br[8] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_11 
+ bl[9] br[9] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_12 
+ bl[10] br[10] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_13 
+ bl[11] br[11] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_14 
+ bl[12] br[12] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_15 
+ bl[13] br[13] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_16 
+ bl[14] br[14] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_17 
+ bl[15] br[15] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_18 
+ bl[16] br[16] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_19 
+ bl[17] br[17] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_20 
+ bl[18] br[18] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_21 
+ bl[19] br[19] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_22 
+ bl[20] br[20] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_23 
+ bl[21] br[21] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_24 
+ bl[22] br[22] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_25 
+ bl[23] br[23] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_26 
+ bl[24] br[24] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_27 
+ bl[25] br[25] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_28 
+ bl[26] br[26] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_29 
+ bl[27] br[27] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_30 
+ bl[28] br[28] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_31 
+ bl[29] br[29] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_32 
+ bl[30] br[30] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_33 
+ bl[31] br[31] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_34 
+ bl[32] br[32] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_35 
+ bl[33] br[33] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_36 
+ bl[34] br[34] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_37 
+ bl[35] br[35] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_38 
+ bl[36] br[36] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_39 
+ bl[37] br[37] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_40 
+ bl[38] br[38] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_41 
+ bl[39] br[39] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_42 
+ bl[40] br[40] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_43 
+ bl[41] br[41] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_44 
+ bl[42] br[42] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_45 
+ bl[43] br[43] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_46 
+ bl[44] br[44] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_47 
+ bl[45] br[45] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_48 
+ bl[46] br[46] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_49 
+ bl[47] br[47] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_50 
+ bl[48] br[48] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_51 
+ bl[49] br[49] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_52 
+ bl[50] br[50] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_53 
+ bl[51] br[51] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_54 
+ bl[52] br[52] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_55 
+ bl[53] br[53] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_56 
+ bl[54] br[54] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_57 
+ bl[55] br[55] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_58 
+ bl[56] br[56] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_59 
+ bl[57] br[57] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_60 
+ bl[58] br[58] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_61 
+ bl[59] br[59] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_62 
+ bl[60] br[60] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_63 
+ bl[61] br[61] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_64 
+ bl[62] br[62] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_65 
+ bl[63] br[63] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_66 
+ bl[64] br[64] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_67 
+ bl[65] br[65] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_68 
+ bl[66] br[66] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_69 
+ bl[67] br[67] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_70 
+ bl[68] br[68] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_71 
+ bl[69] br[69] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_72 
+ bl[70] br[70] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_73 
+ bl[71] br[71] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_74 
+ bl[72] br[72] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_75 
+ bl[73] br[73] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_76 
+ bl[74] br[74] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_77 
+ bl[75] br[75] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_78 
+ bl[76] br[76] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_79 
+ bl[77] br[77] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_80 
+ bl[78] br[78] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_81 
+ bl[79] br[79] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_82 
+ bl[80] br[80] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_83 
+ bl[81] br[81] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_84 
+ bl[82] br[82] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_85 
+ bl[83] br[83] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_86 
+ bl[84] br[84] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_87 
+ bl[85] br[85] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_88 
+ bl[86] br[86] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_89 
+ bl[87] br[87] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_90 
+ bl[88] br[88] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_91 
+ bl[89] br[89] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_92 
+ bl[90] br[90] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_93 
+ bl[91] br[91] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_94 
+ bl[92] br[92] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_95 
+ bl[93] br[93] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_96 
+ bl[94] br[94] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_97 
+ bl[95] br[95] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_98 
+ bl[96] br[96] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_99 
+ bl[97] br[97] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_100 
+ bl[98] br[98] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_101 
+ bl[99] br[99] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_102 
+ bl[100] br[100] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_103 
+ bl[101] br[101] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_104 
+ bl[102] br[102] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_105 
+ bl[103] br[103] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_106 
+ bl[104] br[104] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_107 
+ bl[105] br[105] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_108 
+ bl[106] br[106] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_109 
+ bl[107] br[107] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_110 
+ bl[108] br[108] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_111 
+ bl[109] br[109] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_112 
+ bl[110] br[110] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_113 
+ bl[111] br[111] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_114 
+ bl[112] br[112] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_115 
+ bl[113] br[113] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_116 
+ bl[114] br[114] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_117 
+ bl[115] br[115] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_118 
+ bl[116] br[116] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_119 
+ bl[117] br[117] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_120 
+ bl[118] br[118] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_121 
+ bl[119] br[119] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_122 
+ bl[120] br[120] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_123 
+ bl[121] br[121] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_124 
+ bl[122] br[122] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_125 
+ bl[123] br[123] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_126 
+ bl[124] br[124] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_127 
+ bl[125] br[125] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_128 
+ bl[126] br[126] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_129 
+ bl[127] br[127] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_130 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_131 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_0 
+ vdd vdd vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_1 
+ rbl rbr vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_2 
+ bl[0] br[0] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_3 
+ bl[1] br[1] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_4 
+ bl[2] br[2] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_5 
+ bl[3] br[3] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_6 
+ bl[4] br[4] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_7 
+ bl[5] br[5] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_8 
+ bl[6] br[6] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_9 
+ bl[7] br[7] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_10 
+ bl[8] br[8] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_11 
+ bl[9] br[9] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_12 
+ bl[10] br[10] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_13 
+ bl[11] br[11] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_14 
+ bl[12] br[12] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_15 
+ bl[13] br[13] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_16 
+ bl[14] br[14] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_17 
+ bl[15] br[15] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_18 
+ bl[16] br[16] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_19 
+ bl[17] br[17] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_20 
+ bl[18] br[18] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_21 
+ bl[19] br[19] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_22 
+ bl[20] br[20] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_23 
+ bl[21] br[21] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_24 
+ bl[22] br[22] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_25 
+ bl[23] br[23] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_26 
+ bl[24] br[24] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_27 
+ bl[25] br[25] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_28 
+ bl[26] br[26] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_29 
+ bl[27] br[27] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_30 
+ bl[28] br[28] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_31 
+ bl[29] br[29] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_32 
+ bl[30] br[30] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_33 
+ bl[31] br[31] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_34 
+ bl[32] br[32] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_35 
+ bl[33] br[33] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_36 
+ bl[34] br[34] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_37 
+ bl[35] br[35] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_38 
+ bl[36] br[36] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_39 
+ bl[37] br[37] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_40 
+ bl[38] br[38] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_41 
+ bl[39] br[39] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_42 
+ bl[40] br[40] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_43 
+ bl[41] br[41] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_44 
+ bl[42] br[42] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_45 
+ bl[43] br[43] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_46 
+ bl[44] br[44] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_47 
+ bl[45] br[45] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_48 
+ bl[46] br[46] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_49 
+ bl[47] br[47] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_50 
+ bl[48] br[48] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_51 
+ bl[49] br[49] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_52 
+ bl[50] br[50] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_53 
+ bl[51] br[51] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_54 
+ bl[52] br[52] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_55 
+ bl[53] br[53] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_56 
+ bl[54] br[54] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_57 
+ bl[55] br[55] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_58 
+ bl[56] br[56] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_59 
+ bl[57] br[57] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_60 
+ bl[58] br[58] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_61 
+ bl[59] br[59] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_62 
+ bl[60] br[60] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_63 
+ bl[61] br[61] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_64 
+ bl[62] br[62] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_65 
+ bl[63] br[63] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_66 
+ bl[64] br[64] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_67 
+ bl[65] br[65] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_68 
+ bl[66] br[66] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_69 
+ bl[67] br[67] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_70 
+ bl[68] br[68] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_71 
+ bl[69] br[69] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_72 
+ bl[70] br[70] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_73 
+ bl[71] br[71] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_74 
+ bl[72] br[72] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_75 
+ bl[73] br[73] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_76 
+ bl[74] br[74] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_77 
+ bl[75] br[75] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_78 
+ bl[76] br[76] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_79 
+ bl[77] br[77] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_80 
+ bl[78] br[78] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_81 
+ bl[79] br[79] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_82 
+ bl[80] br[80] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_83 
+ bl[81] br[81] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_84 
+ bl[82] br[82] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_85 
+ bl[83] br[83] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_86 
+ bl[84] br[84] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_87 
+ bl[85] br[85] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_88 
+ bl[86] br[86] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_89 
+ bl[87] br[87] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_90 
+ bl[88] br[88] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_91 
+ bl[89] br[89] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_92 
+ bl[90] br[90] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_93 
+ bl[91] br[91] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_94 
+ bl[92] br[92] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_95 
+ bl[93] br[93] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_96 
+ bl[94] br[94] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_97 
+ bl[95] br[95] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_98 
+ bl[96] br[96] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_99 
+ bl[97] br[97] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_100 
+ bl[98] br[98] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_101 
+ bl[99] br[99] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_102 
+ bl[100] br[100] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_103 
+ bl[101] br[101] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_104 
+ bl[102] br[102] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_105 
+ bl[103] br[103] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_106 
+ bl[104] br[104] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_107 
+ bl[105] br[105] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_108 
+ bl[106] br[106] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_109 
+ bl[107] br[107] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_110 
+ bl[108] br[108] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_111 
+ bl[109] br[109] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_112 
+ bl[110] br[110] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_113 
+ bl[111] br[111] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_114 
+ bl[112] br[112] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_115 
+ bl[113] br[113] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_116 
+ bl[114] br[114] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_117 
+ bl[115] br[115] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_118 
+ bl[116] br[116] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_119 
+ bl[117] br[117] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_120 
+ bl[118] br[118] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_121 
+ bl[119] br[119] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_122 
+ bl[120] br[120] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_123 
+ bl[121] br[121] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_124 
+ bl[122] br[122] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_125 
+ bl[123] br[123] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_126 
+ bl[124] br[124] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_127 
+ bl[125] br[125] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_128 
+ bl[126] br[126] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_129 
+ bl[127] br[127] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_130 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_131 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_0 
+ vdd vdd vss vdd vpb vnb wl[4] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_6_1 
+ rbl rbr vss vdd vpb vnb wl[4] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_6_2 
+ bl[0] br[0] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_3 
+ bl[1] br[1] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_4 
+ bl[2] br[2] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_5 
+ bl[3] br[3] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_6 
+ bl[4] br[4] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_7 
+ bl[5] br[5] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_8 
+ bl[6] br[6] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_9 
+ bl[7] br[7] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_10 
+ bl[8] br[8] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_11 
+ bl[9] br[9] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_12 
+ bl[10] br[10] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_13 
+ bl[11] br[11] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_14 
+ bl[12] br[12] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_15 
+ bl[13] br[13] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_16 
+ bl[14] br[14] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_17 
+ bl[15] br[15] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_18 
+ bl[16] br[16] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_19 
+ bl[17] br[17] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_20 
+ bl[18] br[18] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_21 
+ bl[19] br[19] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_22 
+ bl[20] br[20] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_23 
+ bl[21] br[21] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_24 
+ bl[22] br[22] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_25 
+ bl[23] br[23] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_26 
+ bl[24] br[24] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_27 
+ bl[25] br[25] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_28 
+ bl[26] br[26] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_29 
+ bl[27] br[27] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_30 
+ bl[28] br[28] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_31 
+ bl[29] br[29] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_32 
+ bl[30] br[30] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_33 
+ bl[31] br[31] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_34 
+ bl[32] br[32] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_35 
+ bl[33] br[33] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_36 
+ bl[34] br[34] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_37 
+ bl[35] br[35] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_38 
+ bl[36] br[36] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_39 
+ bl[37] br[37] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_40 
+ bl[38] br[38] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_41 
+ bl[39] br[39] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_42 
+ bl[40] br[40] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_43 
+ bl[41] br[41] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_44 
+ bl[42] br[42] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_45 
+ bl[43] br[43] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_46 
+ bl[44] br[44] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_47 
+ bl[45] br[45] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_48 
+ bl[46] br[46] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_49 
+ bl[47] br[47] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_50 
+ bl[48] br[48] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_51 
+ bl[49] br[49] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_52 
+ bl[50] br[50] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_53 
+ bl[51] br[51] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_54 
+ bl[52] br[52] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_55 
+ bl[53] br[53] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_56 
+ bl[54] br[54] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_57 
+ bl[55] br[55] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_58 
+ bl[56] br[56] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_59 
+ bl[57] br[57] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_60 
+ bl[58] br[58] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_61 
+ bl[59] br[59] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_62 
+ bl[60] br[60] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_63 
+ bl[61] br[61] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_64 
+ bl[62] br[62] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_65 
+ bl[63] br[63] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_66 
+ bl[64] br[64] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_67 
+ bl[65] br[65] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_68 
+ bl[66] br[66] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_69 
+ bl[67] br[67] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_70 
+ bl[68] br[68] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_71 
+ bl[69] br[69] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_72 
+ bl[70] br[70] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_73 
+ bl[71] br[71] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_74 
+ bl[72] br[72] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_75 
+ bl[73] br[73] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_76 
+ bl[74] br[74] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_77 
+ bl[75] br[75] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_78 
+ bl[76] br[76] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_79 
+ bl[77] br[77] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_80 
+ bl[78] br[78] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_81 
+ bl[79] br[79] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_82 
+ bl[80] br[80] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_83 
+ bl[81] br[81] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_84 
+ bl[82] br[82] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_85 
+ bl[83] br[83] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_86 
+ bl[84] br[84] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_87 
+ bl[85] br[85] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_88 
+ bl[86] br[86] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_89 
+ bl[87] br[87] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_90 
+ bl[88] br[88] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_91 
+ bl[89] br[89] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_92 
+ bl[90] br[90] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_93 
+ bl[91] br[91] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_94 
+ bl[92] br[92] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_95 
+ bl[93] br[93] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_96 
+ bl[94] br[94] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_97 
+ bl[95] br[95] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_98 
+ bl[96] br[96] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_99 
+ bl[97] br[97] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_100 
+ bl[98] br[98] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_101 
+ bl[99] br[99] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_102 
+ bl[100] br[100] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_103 
+ bl[101] br[101] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_104 
+ bl[102] br[102] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_105 
+ bl[103] br[103] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_106 
+ bl[104] br[104] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_107 
+ bl[105] br[105] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_108 
+ bl[106] br[106] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_109 
+ bl[107] br[107] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_110 
+ bl[108] br[108] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_111 
+ bl[109] br[109] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_112 
+ bl[110] br[110] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_113 
+ bl[111] br[111] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_114 
+ bl[112] br[112] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_115 
+ bl[113] br[113] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_116 
+ bl[114] br[114] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_117 
+ bl[115] br[115] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_118 
+ bl[116] br[116] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_119 
+ bl[117] br[117] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_120 
+ bl[118] br[118] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_121 
+ bl[119] br[119] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_122 
+ bl[120] br[120] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_123 
+ bl[121] br[121] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_124 
+ bl[122] br[122] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_125 
+ bl[123] br[123] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_126 
+ bl[124] br[124] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_127 
+ bl[125] br[125] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_128 
+ bl[126] br[126] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_129 
+ bl[127] br[127] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_130 
+ vdd vdd vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_131 
+ vdd vdd vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_0 
+ vdd vdd vss vdd vpb vnb wl[5] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_7_1 
+ rbl rbr vss vdd vpb vnb wl[5] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_7_2 
+ bl[0] br[0] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_3 
+ bl[1] br[1] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_4 
+ bl[2] br[2] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_5 
+ bl[3] br[3] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_6 
+ bl[4] br[4] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_7 
+ bl[5] br[5] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_8 
+ bl[6] br[6] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_9 
+ bl[7] br[7] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_10 
+ bl[8] br[8] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_11 
+ bl[9] br[9] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_12 
+ bl[10] br[10] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_13 
+ bl[11] br[11] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_14 
+ bl[12] br[12] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_15 
+ bl[13] br[13] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_16 
+ bl[14] br[14] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_17 
+ bl[15] br[15] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_18 
+ bl[16] br[16] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_19 
+ bl[17] br[17] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_20 
+ bl[18] br[18] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_21 
+ bl[19] br[19] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_22 
+ bl[20] br[20] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_23 
+ bl[21] br[21] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_24 
+ bl[22] br[22] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_25 
+ bl[23] br[23] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_26 
+ bl[24] br[24] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_27 
+ bl[25] br[25] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_28 
+ bl[26] br[26] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_29 
+ bl[27] br[27] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_30 
+ bl[28] br[28] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_31 
+ bl[29] br[29] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_32 
+ bl[30] br[30] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_33 
+ bl[31] br[31] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_34 
+ bl[32] br[32] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_35 
+ bl[33] br[33] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_36 
+ bl[34] br[34] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_37 
+ bl[35] br[35] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_38 
+ bl[36] br[36] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_39 
+ bl[37] br[37] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_40 
+ bl[38] br[38] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_41 
+ bl[39] br[39] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_42 
+ bl[40] br[40] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_43 
+ bl[41] br[41] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_44 
+ bl[42] br[42] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_45 
+ bl[43] br[43] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_46 
+ bl[44] br[44] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_47 
+ bl[45] br[45] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_48 
+ bl[46] br[46] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_49 
+ bl[47] br[47] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_50 
+ bl[48] br[48] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_51 
+ bl[49] br[49] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_52 
+ bl[50] br[50] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_53 
+ bl[51] br[51] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_54 
+ bl[52] br[52] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_55 
+ bl[53] br[53] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_56 
+ bl[54] br[54] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_57 
+ bl[55] br[55] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_58 
+ bl[56] br[56] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_59 
+ bl[57] br[57] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_60 
+ bl[58] br[58] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_61 
+ bl[59] br[59] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_62 
+ bl[60] br[60] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_63 
+ bl[61] br[61] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_64 
+ bl[62] br[62] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_65 
+ bl[63] br[63] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_66 
+ bl[64] br[64] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_67 
+ bl[65] br[65] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_68 
+ bl[66] br[66] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_69 
+ bl[67] br[67] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_70 
+ bl[68] br[68] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_71 
+ bl[69] br[69] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_72 
+ bl[70] br[70] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_73 
+ bl[71] br[71] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_74 
+ bl[72] br[72] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_75 
+ bl[73] br[73] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_76 
+ bl[74] br[74] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_77 
+ bl[75] br[75] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_78 
+ bl[76] br[76] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_79 
+ bl[77] br[77] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_80 
+ bl[78] br[78] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_81 
+ bl[79] br[79] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_82 
+ bl[80] br[80] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_83 
+ bl[81] br[81] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_84 
+ bl[82] br[82] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_85 
+ bl[83] br[83] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_86 
+ bl[84] br[84] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_87 
+ bl[85] br[85] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_88 
+ bl[86] br[86] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_89 
+ bl[87] br[87] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_90 
+ bl[88] br[88] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_91 
+ bl[89] br[89] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_92 
+ bl[90] br[90] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_93 
+ bl[91] br[91] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_94 
+ bl[92] br[92] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_95 
+ bl[93] br[93] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_96 
+ bl[94] br[94] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_97 
+ bl[95] br[95] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_98 
+ bl[96] br[96] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_99 
+ bl[97] br[97] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_100 
+ bl[98] br[98] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_101 
+ bl[99] br[99] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_102 
+ bl[100] br[100] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_103 
+ bl[101] br[101] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_104 
+ bl[102] br[102] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_105 
+ bl[103] br[103] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_106 
+ bl[104] br[104] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_107 
+ bl[105] br[105] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_108 
+ bl[106] br[106] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_109 
+ bl[107] br[107] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_110 
+ bl[108] br[108] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_111 
+ bl[109] br[109] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_112 
+ bl[110] br[110] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_113 
+ bl[111] br[111] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_114 
+ bl[112] br[112] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_115 
+ bl[113] br[113] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_116 
+ bl[114] br[114] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_117 
+ bl[115] br[115] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_118 
+ bl[116] br[116] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_119 
+ bl[117] br[117] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_120 
+ bl[118] br[118] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_121 
+ bl[119] br[119] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_122 
+ bl[120] br[120] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_123 
+ bl[121] br[121] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_124 
+ bl[122] br[122] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_125 
+ bl[123] br[123] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_126 
+ bl[124] br[124] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_127 
+ bl[125] br[125] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_128 
+ bl[126] br[126] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_129 
+ bl[127] br[127] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_130 
+ vdd vdd vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_131 
+ vdd vdd vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_0 
+ vdd vdd vss vdd vpb vnb wl[6] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_8_1 
+ rbl rbr vss vdd vpb vnb wl[6] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_8_2 
+ bl[0] br[0] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_3 
+ bl[1] br[1] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_4 
+ bl[2] br[2] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_5 
+ bl[3] br[3] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_6 
+ bl[4] br[4] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_7 
+ bl[5] br[5] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_8 
+ bl[6] br[6] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_9 
+ bl[7] br[7] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_10 
+ bl[8] br[8] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_11 
+ bl[9] br[9] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_12 
+ bl[10] br[10] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_13 
+ bl[11] br[11] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_14 
+ bl[12] br[12] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_15 
+ bl[13] br[13] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_16 
+ bl[14] br[14] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_17 
+ bl[15] br[15] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_18 
+ bl[16] br[16] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_19 
+ bl[17] br[17] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_20 
+ bl[18] br[18] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_21 
+ bl[19] br[19] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_22 
+ bl[20] br[20] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_23 
+ bl[21] br[21] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_24 
+ bl[22] br[22] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_25 
+ bl[23] br[23] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_26 
+ bl[24] br[24] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_27 
+ bl[25] br[25] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_28 
+ bl[26] br[26] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_29 
+ bl[27] br[27] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_30 
+ bl[28] br[28] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_31 
+ bl[29] br[29] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_32 
+ bl[30] br[30] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_33 
+ bl[31] br[31] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_34 
+ bl[32] br[32] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_35 
+ bl[33] br[33] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_36 
+ bl[34] br[34] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_37 
+ bl[35] br[35] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_38 
+ bl[36] br[36] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_39 
+ bl[37] br[37] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_40 
+ bl[38] br[38] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_41 
+ bl[39] br[39] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_42 
+ bl[40] br[40] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_43 
+ bl[41] br[41] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_44 
+ bl[42] br[42] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_45 
+ bl[43] br[43] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_46 
+ bl[44] br[44] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_47 
+ bl[45] br[45] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_48 
+ bl[46] br[46] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_49 
+ bl[47] br[47] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_50 
+ bl[48] br[48] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_51 
+ bl[49] br[49] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_52 
+ bl[50] br[50] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_53 
+ bl[51] br[51] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_54 
+ bl[52] br[52] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_55 
+ bl[53] br[53] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_56 
+ bl[54] br[54] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_57 
+ bl[55] br[55] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_58 
+ bl[56] br[56] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_59 
+ bl[57] br[57] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_60 
+ bl[58] br[58] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_61 
+ bl[59] br[59] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_62 
+ bl[60] br[60] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_63 
+ bl[61] br[61] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_64 
+ bl[62] br[62] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_65 
+ bl[63] br[63] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_66 
+ bl[64] br[64] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_67 
+ bl[65] br[65] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_68 
+ bl[66] br[66] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_69 
+ bl[67] br[67] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_70 
+ bl[68] br[68] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_71 
+ bl[69] br[69] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_72 
+ bl[70] br[70] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_73 
+ bl[71] br[71] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_74 
+ bl[72] br[72] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_75 
+ bl[73] br[73] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_76 
+ bl[74] br[74] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_77 
+ bl[75] br[75] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_78 
+ bl[76] br[76] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_79 
+ bl[77] br[77] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_80 
+ bl[78] br[78] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_81 
+ bl[79] br[79] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_82 
+ bl[80] br[80] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_83 
+ bl[81] br[81] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_84 
+ bl[82] br[82] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_85 
+ bl[83] br[83] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_86 
+ bl[84] br[84] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_87 
+ bl[85] br[85] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_88 
+ bl[86] br[86] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_89 
+ bl[87] br[87] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_90 
+ bl[88] br[88] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_91 
+ bl[89] br[89] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_92 
+ bl[90] br[90] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_93 
+ bl[91] br[91] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_94 
+ bl[92] br[92] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_95 
+ bl[93] br[93] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_96 
+ bl[94] br[94] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_97 
+ bl[95] br[95] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_98 
+ bl[96] br[96] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_99 
+ bl[97] br[97] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_100 
+ bl[98] br[98] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_101 
+ bl[99] br[99] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_102 
+ bl[100] br[100] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_103 
+ bl[101] br[101] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_104 
+ bl[102] br[102] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_105 
+ bl[103] br[103] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_106 
+ bl[104] br[104] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_107 
+ bl[105] br[105] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_108 
+ bl[106] br[106] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_109 
+ bl[107] br[107] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_110 
+ bl[108] br[108] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_111 
+ bl[109] br[109] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_112 
+ bl[110] br[110] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_113 
+ bl[111] br[111] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_114 
+ bl[112] br[112] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_115 
+ bl[113] br[113] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_116 
+ bl[114] br[114] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_117 
+ bl[115] br[115] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_118 
+ bl[116] br[116] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_119 
+ bl[117] br[117] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_120 
+ bl[118] br[118] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_121 
+ bl[119] br[119] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_122 
+ bl[120] br[120] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_123 
+ bl[121] br[121] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_124 
+ bl[122] br[122] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_125 
+ bl[123] br[123] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_126 
+ bl[124] br[124] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_127 
+ bl[125] br[125] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_128 
+ bl[126] br[126] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_129 
+ bl[127] br[127] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_130 
+ vdd vdd vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_131 
+ vdd vdd vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_0 
+ vdd vdd vss vdd vpb vnb wl[7] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_9_1 
+ rbl rbr vss vdd vpb vnb wl[7] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_9_2 
+ bl[0] br[0] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_3 
+ bl[1] br[1] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_4 
+ bl[2] br[2] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_5 
+ bl[3] br[3] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_6 
+ bl[4] br[4] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_7 
+ bl[5] br[5] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_8 
+ bl[6] br[6] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_9 
+ bl[7] br[7] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_10 
+ bl[8] br[8] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_11 
+ bl[9] br[9] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_12 
+ bl[10] br[10] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_13 
+ bl[11] br[11] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_14 
+ bl[12] br[12] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_15 
+ bl[13] br[13] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_16 
+ bl[14] br[14] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_17 
+ bl[15] br[15] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_18 
+ bl[16] br[16] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_19 
+ bl[17] br[17] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_20 
+ bl[18] br[18] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_21 
+ bl[19] br[19] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_22 
+ bl[20] br[20] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_23 
+ bl[21] br[21] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_24 
+ bl[22] br[22] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_25 
+ bl[23] br[23] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_26 
+ bl[24] br[24] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_27 
+ bl[25] br[25] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_28 
+ bl[26] br[26] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_29 
+ bl[27] br[27] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_30 
+ bl[28] br[28] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_31 
+ bl[29] br[29] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_32 
+ bl[30] br[30] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_33 
+ bl[31] br[31] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_34 
+ bl[32] br[32] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_35 
+ bl[33] br[33] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_36 
+ bl[34] br[34] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_37 
+ bl[35] br[35] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_38 
+ bl[36] br[36] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_39 
+ bl[37] br[37] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_40 
+ bl[38] br[38] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_41 
+ bl[39] br[39] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_42 
+ bl[40] br[40] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_43 
+ bl[41] br[41] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_44 
+ bl[42] br[42] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_45 
+ bl[43] br[43] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_46 
+ bl[44] br[44] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_47 
+ bl[45] br[45] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_48 
+ bl[46] br[46] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_49 
+ bl[47] br[47] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_50 
+ bl[48] br[48] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_51 
+ bl[49] br[49] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_52 
+ bl[50] br[50] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_53 
+ bl[51] br[51] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_54 
+ bl[52] br[52] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_55 
+ bl[53] br[53] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_56 
+ bl[54] br[54] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_57 
+ bl[55] br[55] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_58 
+ bl[56] br[56] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_59 
+ bl[57] br[57] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_60 
+ bl[58] br[58] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_61 
+ bl[59] br[59] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_62 
+ bl[60] br[60] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_63 
+ bl[61] br[61] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_64 
+ bl[62] br[62] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_65 
+ bl[63] br[63] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_66 
+ bl[64] br[64] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_67 
+ bl[65] br[65] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_68 
+ bl[66] br[66] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_69 
+ bl[67] br[67] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_70 
+ bl[68] br[68] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_71 
+ bl[69] br[69] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_72 
+ bl[70] br[70] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_73 
+ bl[71] br[71] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_74 
+ bl[72] br[72] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_75 
+ bl[73] br[73] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_76 
+ bl[74] br[74] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_77 
+ bl[75] br[75] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_78 
+ bl[76] br[76] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_79 
+ bl[77] br[77] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_80 
+ bl[78] br[78] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_81 
+ bl[79] br[79] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_82 
+ bl[80] br[80] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_83 
+ bl[81] br[81] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_84 
+ bl[82] br[82] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_85 
+ bl[83] br[83] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_86 
+ bl[84] br[84] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_87 
+ bl[85] br[85] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_88 
+ bl[86] br[86] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_89 
+ bl[87] br[87] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_90 
+ bl[88] br[88] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_91 
+ bl[89] br[89] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_92 
+ bl[90] br[90] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_93 
+ bl[91] br[91] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_94 
+ bl[92] br[92] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_95 
+ bl[93] br[93] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_96 
+ bl[94] br[94] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_97 
+ bl[95] br[95] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_98 
+ bl[96] br[96] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_99 
+ bl[97] br[97] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_100 
+ bl[98] br[98] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_101 
+ bl[99] br[99] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_102 
+ bl[100] br[100] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_103 
+ bl[101] br[101] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_104 
+ bl[102] br[102] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_105 
+ bl[103] br[103] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_106 
+ bl[104] br[104] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_107 
+ bl[105] br[105] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_108 
+ bl[106] br[106] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_109 
+ bl[107] br[107] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_110 
+ bl[108] br[108] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_111 
+ bl[109] br[109] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_112 
+ bl[110] br[110] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_113 
+ bl[111] br[111] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_114 
+ bl[112] br[112] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_115 
+ bl[113] br[113] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_116 
+ bl[114] br[114] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_117 
+ bl[115] br[115] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_118 
+ bl[116] br[116] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_119 
+ bl[117] br[117] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_120 
+ bl[118] br[118] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_121 
+ bl[119] br[119] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_122 
+ bl[120] br[120] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_123 
+ bl[121] br[121] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_124 
+ bl[122] br[122] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_125 
+ bl[123] br[123] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_126 
+ bl[124] br[124] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_127 
+ bl[125] br[125] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_128 
+ bl[126] br[126] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_129 
+ bl[127] br[127] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_130 
+ vdd vdd vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_131 
+ vdd vdd vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_0 
+ vdd vdd vss vdd vpb vnb wl[8] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_10_1 
+ rbl rbr vss vdd vpb vnb wl[8] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_10_2 
+ bl[0] br[0] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_3 
+ bl[1] br[1] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_4 
+ bl[2] br[2] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_5 
+ bl[3] br[3] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_6 
+ bl[4] br[4] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_7 
+ bl[5] br[5] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_8 
+ bl[6] br[6] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_9 
+ bl[7] br[7] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_10 
+ bl[8] br[8] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_11 
+ bl[9] br[9] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_12 
+ bl[10] br[10] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_13 
+ bl[11] br[11] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_14 
+ bl[12] br[12] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_15 
+ bl[13] br[13] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_16 
+ bl[14] br[14] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_17 
+ bl[15] br[15] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_18 
+ bl[16] br[16] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_19 
+ bl[17] br[17] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_20 
+ bl[18] br[18] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_21 
+ bl[19] br[19] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_22 
+ bl[20] br[20] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_23 
+ bl[21] br[21] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_24 
+ bl[22] br[22] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_25 
+ bl[23] br[23] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_26 
+ bl[24] br[24] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_27 
+ bl[25] br[25] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_28 
+ bl[26] br[26] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_29 
+ bl[27] br[27] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_30 
+ bl[28] br[28] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_31 
+ bl[29] br[29] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_32 
+ bl[30] br[30] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_33 
+ bl[31] br[31] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_34 
+ bl[32] br[32] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_35 
+ bl[33] br[33] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_36 
+ bl[34] br[34] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_37 
+ bl[35] br[35] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_38 
+ bl[36] br[36] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_39 
+ bl[37] br[37] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_40 
+ bl[38] br[38] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_41 
+ bl[39] br[39] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_42 
+ bl[40] br[40] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_43 
+ bl[41] br[41] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_44 
+ bl[42] br[42] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_45 
+ bl[43] br[43] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_46 
+ bl[44] br[44] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_47 
+ bl[45] br[45] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_48 
+ bl[46] br[46] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_49 
+ bl[47] br[47] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_50 
+ bl[48] br[48] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_51 
+ bl[49] br[49] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_52 
+ bl[50] br[50] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_53 
+ bl[51] br[51] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_54 
+ bl[52] br[52] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_55 
+ bl[53] br[53] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_56 
+ bl[54] br[54] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_57 
+ bl[55] br[55] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_58 
+ bl[56] br[56] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_59 
+ bl[57] br[57] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_60 
+ bl[58] br[58] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_61 
+ bl[59] br[59] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_62 
+ bl[60] br[60] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_63 
+ bl[61] br[61] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_64 
+ bl[62] br[62] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_65 
+ bl[63] br[63] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_66 
+ bl[64] br[64] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_67 
+ bl[65] br[65] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_68 
+ bl[66] br[66] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_69 
+ bl[67] br[67] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_70 
+ bl[68] br[68] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_71 
+ bl[69] br[69] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_72 
+ bl[70] br[70] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_73 
+ bl[71] br[71] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_74 
+ bl[72] br[72] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_75 
+ bl[73] br[73] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_76 
+ bl[74] br[74] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_77 
+ bl[75] br[75] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_78 
+ bl[76] br[76] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_79 
+ bl[77] br[77] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_80 
+ bl[78] br[78] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_81 
+ bl[79] br[79] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_82 
+ bl[80] br[80] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_83 
+ bl[81] br[81] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_84 
+ bl[82] br[82] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_85 
+ bl[83] br[83] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_86 
+ bl[84] br[84] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_87 
+ bl[85] br[85] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_88 
+ bl[86] br[86] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_89 
+ bl[87] br[87] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_90 
+ bl[88] br[88] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_91 
+ bl[89] br[89] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_92 
+ bl[90] br[90] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_93 
+ bl[91] br[91] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_94 
+ bl[92] br[92] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_95 
+ bl[93] br[93] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_96 
+ bl[94] br[94] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_97 
+ bl[95] br[95] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_98 
+ bl[96] br[96] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_99 
+ bl[97] br[97] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_100 
+ bl[98] br[98] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_101 
+ bl[99] br[99] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_102 
+ bl[100] br[100] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_103 
+ bl[101] br[101] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_104 
+ bl[102] br[102] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_105 
+ bl[103] br[103] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_106 
+ bl[104] br[104] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_107 
+ bl[105] br[105] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_108 
+ bl[106] br[106] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_109 
+ bl[107] br[107] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_110 
+ bl[108] br[108] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_111 
+ bl[109] br[109] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_112 
+ bl[110] br[110] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_113 
+ bl[111] br[111] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_114 
+ bl[112] br[112] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_115 
+ bl[113] br[113] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_116 
+ bl[114] br[114] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_117 
+ bl[115] br[115] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_118 
+ bl[116] br[116] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_119 
+ bl[117] br[117] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_120 
+ bl[118] br[118] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_121 
+ bl[119] br[119] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_122 
+ bl[120] br[120] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_123 
+ bl[121] br[121] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_124 
+ bl[122] br[122] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_125 
+ bl[123] br[123] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_126 
+ bl[124] br[124] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_127 
+ bl[125] br[125] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_128 
+ bl[126] br[126] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_129 
+ bl[127] br[127] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_130 
+ vdd vdd vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_131 
+ vdd vdd vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_0 
+ vdd vdd vss vdd vpb vnb wl[9] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_11_1 
+ rbl rbr vss vdd vpb vnb wl[9] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_11_2 
+ bl[0] br[0] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_3 
+ bl[1] br[1] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_4 
+ bl[2] br[2] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_5 
+ bl[3] br[3] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_6 
+ bl[4] br[4] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_7 
+ bl[5] br[5] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_8 
+ bl[6] br[6] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_9 
+ bl[7] br[7] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_10 
+ bl[8] br[8] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_11 
+ bl[9] br[9] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_12 
+ bl[10] br[10] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_13 
+ bl[11] br[11] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_14 
+ bl[12] br[12] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_15 
+ bl[13] br[13] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_16 
+ bl[14] br[14] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_17 
+ bl[15] br[15] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_18 
+ bl[16] br[16] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_19 
+ bl[17] br[17] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_20 
+ bl[18] br[18] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_21 
+ bl[19] br[19] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_22 
+ bl[20] br[20] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_23 
+ bl[21] br[21] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_24 
+ bl[22] br[22] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_25 
+ bl[23] br[23] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_26 
+ bl[24] br[24] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_27 
+ bl[25] br[25] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_28 
+ bl[26] br[26] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_29 
+ bl[27] br[27] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_30 
+ bl[28] br[28] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_31 
+ bl[29] br[29] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_32 
+ bl[30] br[30] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_33 
+ bl[31] br[31] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_34 
+ bl[32] br[32] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_35 
+ bl[33] br[33] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_36 
+ bl[34] br[34] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_37 
+ bl[35] br[35] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_38 
+ bl[36] br[36] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_39 
+ bl[37] br[37] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_40 
+ bl[38] br[38] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_41 
+ bl[39] br[39] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_42 
+ bl[40] br[40] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_43 
+ bl[41] br[41] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_44 
+ bl[42] br[42] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_45 
+ bl[43] br[43] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_46 
+ bl[44] br[44] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_47 
+ bl[45] br[45] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_48 
+ bl[46] br[46] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_49 
+ bl[47] br[47] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_50 
+ bl[48] br[48] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_51 
+ bl[49] br[49] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_52 
+ bl[50] br[50] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_53 
+ bl[51] br[51] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_54 
+ bl[52] br[52] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_55 
+ bl[53] br[53] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_56 
+ bl[54] br[54] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_57 
+ bl[55] br[55] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_58 
+ bl[56] br[56] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_59 
+ bl[57] br[57] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_60 
+ bl[58] br[58] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_61 
+ bl[59] br[59] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_62 
+ bl[60] br[60] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_63 
+ bl[61] br[61] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_64 
+ bl[62] br[62] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_65 
+ bl[63] br[63] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_66 
+ bl[64] br[64] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_67 
+ bl[65] br[65] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_68 
+ bl[66] br[66] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_69 
+ bl[67] br[67] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_70 
+ bl[68] br[68] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_71 
+ bl[69] br[69] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_72 
+ bl[70] br[70] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_73 
+ bl[71] br[71] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_74 
+ bl[72] br[72] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_75 
+ bl[73] br[73] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_76 
+ bl[74] br[74] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_77 
+ bl[75] br[75] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_78 
+ bl[76] br[76] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_79 
+ bl[77] br[77] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_80 
+ bl[78] br[78] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_81 
+ bl[79] br[79] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_82 
+ bl[80] br[80] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_83 
+ bl[81] br[81] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_84 
+ bl[82] br[82] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_85 
+ bl[83] br[83] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_86 
+ bl[84] br[84] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_87 
+ bl[85] br[85] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_88 
+ bl[86] br[86] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_89 
+ bl[87] br[87] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_90 
+ bl[88] br[88] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_91 
+ bl[89] br[89] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_92 
+ bl[90] br[90] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_93 
+ bl[91] br[91] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_94 
+ bl[92] br[92] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_95 
+ bl[93] br[93] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_96 
+ bl[94] br[94] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_97 
+ bl[95] br[95] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_98 
+ bl[96] br[96] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_99 
+ bl[97] br[97] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_100 
+ bl[98] br[98] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_101 
+ bl[99] br[99] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_102 
+ bl[100] br[100] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_103 
+ bl[101] br[101] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_104 
+ bl[102] br[102] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_105 
+ bl[103] br[103] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_106 
+ bl[104] br[104] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_107 
+ bl[105] br[105] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_108 
+ bl[106] br[106] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_109 
+ bl[107] br[107] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_110 
+ bl[108] br[108] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_111 
+ bl[109] br[109] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_112 
+ bl[110] br[110] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_113 
+ bl[111] br[111] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_114 
+ bl[112] br[112] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_115 
+ bl[113] br[113] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_116 
+ bl[114] br[114] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_117 
+ bl[115] br[115] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_118 
+ bl[116] br[116] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_119 
+ bl[117] br[117] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_120 
+ bl[118] br[118] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_121 
+ bl[119] br[119] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_122 
+ bl[120] br[120] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_123 
+ bl[121] br[121] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_124 
+ bl[122] br[122] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_125 
+ bl[123] br[123] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_126 
+ bl[124] br[124] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_127 
+ bl[125] br[125] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_128 
+ bl[126] br[126] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_129 
+ bl[127] br[127] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_130 
+ vdd vdd vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_131 
+ vdd vdd vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_0 
+ vdd vdd vss vdd vpb vnb wl[10] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_12_1 
+ rbl rbr vss vdd vpb vnb wl[10] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_12_2 
+ bl[0] br[0] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_3 
+ bl[1] br[1] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_4 
+ bl[2] br[2] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_5 
+ bl[3] br[3] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_6 
+ bl[4] br[4] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_7 
+ bl[5] br[5] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_8 
+ bl[6] br[6] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_9 
+ bl[7] br[7] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_10 
+ bl[8] br[8] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_11 
+ bl[9] br[9] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_12 
+ bl[10] br[10] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_13 
+ bl[11] br[11] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_14 
+ bl[12] br[12] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_15 
+ bl[13] br[13] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_16 
+ bl[14] br[14] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_17 
+ bl[15] br[15] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_18 
+ bl[16] br[16] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_19 
+ bl[17] br[17] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_20 
+ bl[18] br[18] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_21 
+ bl[19] br[19] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_22 
+ bl[20] br[20] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_23 
+ bl[21] br[21] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_24 
+ bl[22] br[22] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_25 
+ bl[23] br[23] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_26 
+ bl[24] br[24] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_27 
+ bl[25] br[25] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_28 
+ bl[26] br[26] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_29 
+ bl[27] br[27] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_30 
+ bl[28] br[28] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_31 
+ bl[29] br[29] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_32 
+ bl[30] br[30] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_33 
+ bl[31] br[31] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_34 
+ bl[32] br[32] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_35 
+ bl[33] br[33] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_36 
+ bl[34] br[34] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_37 
+ bl[35] br[35] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_38 
+ bl[36] br[36] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_39 
+ bl[37] br[37] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_40 
+ bl[38] br[38] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_41 
+ bl[39] br[39] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_42 
+ bl[40] br[40] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_43 
+ bl[41] br[41] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_44 
+ bl[42] br[42] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_45 
+ bl[43] br[43] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_46 
+ bl[44] br[44] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_47 
+ bl[45] br[45] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_48 
+ bl[46] br[46] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_49 
+ bl[47] br[47] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_50 
+ bl[48] br[48] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_51 
+ bl[49] br[49] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_52 
+ bl[50] br[50] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_53 
+ bl[51] br[51] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_54 
+ bl[52] br[52] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_55 
+ bl[53] br[53] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_56 
+ bl[54] br[54] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_57 
+ bl[55] br[55] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_58 
+ bl[56] br[56] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_59 
+ bl[57] br[57] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_60 
+ bl[58] br[58] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_61 
+ bl[59] br[59] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_62 
+ bl[60] br[60] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_63 
+ bl[61] br[61] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_64 
+ bl[62] br[62] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_65 
+ bl[63] br[63] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_66 
+ bl[64] br[64] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_67 
+ bl[65] br[65] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_68 
+ bl[66] br[66] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_69 
+ bl[67] br[67] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_70 
+ bl[68] br[68] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_71 
+ bl[69] br[69] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_72 
+ bl[70] br[70] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_73 
+ bl[71] br[71] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_74 
+ bl[72] br[72] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_75 
+ bl[73] br[73] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_76 
+ bl[74] br[74] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_77 
+ bl[75] br[75] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_78 
+ bl[76] br[76] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_79 
+ bl[77] br[77] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_80 
+ bl[78] br[78] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_81 
+ bl[79] br[79] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_82 
+ bl[80] br[80] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_83 
+ bl[81] br[81] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_84 
+ bl[82] br[82] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_85 
+ bl[83] br[83] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_86 
+ bl[84] br[84] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_87 
+ bl[85] br[85] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_88 
+ bl[86] br[86] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_89 
+ bl[87] br[87] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_90 
+ bl[88] br[88] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_91 
+ bl[89] br[89] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_92 
+ bl[90] br[90] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_93 
+ bl[91] br[91] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_94 
+ bl[92] br[92] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_95 
+ bl[93] br[93] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_96 
+ bl[94] br[94] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_97 
+ bl[95] br[95] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_98 
+ bl[96] br[96] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_99 
+ bl[97] br[97] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_100 
+ bl[98] br[98] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_101 
+ bl[99] br[99] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_102 
+ bl[100] br[100] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_103 
+ bl[101] br[101] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_104 
+ bl[102] br[102] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_105 
+ bl[103] br[103] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_106 
+ bl[104] br[104] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_107 
+ bl[105] br[105] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_108 
+ bl[106] br[106] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_109 
+ bl[107] br[107] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_110 
+ bl[108] br[108] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_111 
+ bl[109] br[109] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_112 
+ bl[110] br[110] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_113 
+ bl[111] br[111] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_114 
+ bl[112] br[112] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_115 
+ bl[113] br[113] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_116 
+ bl[114] br[114] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_117 
+ bl[115] br[115] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_118 
+ bl[116] br[116] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_119 
+ bl[117] br[117] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_120 
+ bl[118] br[118] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_121 
+ bl[119] br[119] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_122 
+ bl[120] br[120] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_123 
+ bl[121] br[121] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_124 
+ bl[122] br[122] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_125 
+ bl[123] br[123] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_126 
+ bl[124] br[124] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_127 
+ bl[125] br[125] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_128 
+ bl[126] br[126] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_129 
+ bl[127] br[127] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_130 
+ vdd vdd vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_131 
+ vdd vdd vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_0 
+ vdd vdd vss vdd vpb vnb wl[11] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_13_1 
+ rbl rbr vss vdd vpb vnb wl[11] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_13_2 
+ bl[0] br[0] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_3 
+ bl[1] br[1] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_4 
+ bl[2] br[2] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_5 
+ bl[3] br[3] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_6 
+ bl[4] br[4] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_7 
+ bl[5] br[5] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_8 
+ bl[6] br[6] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_9 
+ bl[7] br[7] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_10 
+ bl[8] br[8] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_11 
+ bl[9] br[9] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_12 
+ bl[10] br[10] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_13 
+ bl[11] br[11] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_14 
+ bl[12] br[12] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_15 
+ bl[13] br[13] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_16 
+ bl[14] br[14] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_17 
+ bl[15] br[15] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_18 
+ bl[16] br[16] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_19 
+ bl[17] br[17] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_20 
+ bl[18] br[18] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_21 
+ bl[19] br[19] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_22 
+ bl[20] br[20] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_23 
+ bl[21] br[21] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_24 
+ bl[22] br[22] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_25 
+ bl[23] br[23] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_26 
+ bl[24] br[24] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_27 
+ bl[25] br[25] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_28 
+ bl[26] br[26] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_29 
+ bl[27] br[27] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_30 
+ bl[28] br[28] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_31 
+ bl[29] br[29] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_32 
+ bl[30] br[30] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_33 
+ bl[31] br[31] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_34 
+ bl[32] br[32] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_35 
+ bl[33] br[33] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_36 
+ bl[34] br[34] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_37 
+ bl[35] br[35] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_38 
+ bl[36] br[36] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_39 
+ bl[37] br[37] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_40 
+ bl[38] br[38] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_41 
+ bl[39] br[39] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_42 
+ bl[40] br[40] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_43 
+ bl[41] br[41] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_44 
+ bl[42] br[42] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_45 
+ bl[43] br[43] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_46 
+ bl[44] br[44] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_47 
+ bl[45] br[45] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_48 
+ bl[46] br[46] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_49 
+ bl[47] br[47] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_50 
+ bl[48] br[48] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_51 
+ bl[49] br[49] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_52 
+ bl[50] br[50] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_53 
+ bl[51] br[51] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_54 
+ bl[52] br[52] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_55 
+ bl[53] br[53] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_56 
+ bl[54] br[54] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_57 
+ bl[55] br[55] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_58 
+ bl[56] br[56] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_59 
+ bl[57] br[57] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_60 
+ bl[58] br[58] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_61 
+ bl[59] br[59] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_62 
+ bl[60] br[60] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_63 
+ bl[61] br[61] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_64 
+ bl[62] br[62] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_65 
+ bl[63] br[63] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_66 
+ bl[64] br[64] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_67 
+ bl[65] br[65] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_68 
+ bl[66] br[66] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_69 
+ bl[67] br[67] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_70 
+ bl[68] br[68] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_71 
+ bl[69] br[69] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_72 
+ bl[70] br[70] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_73 
+ bl[71] br[71] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_74 
+ bl[72] br[72] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_75 
+ bl[73] br[73] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_76 
+ bl[74] br[74] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_77 
+ bl[75] br[75] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_78 
+ bl[76] br[76] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_79 
+ bl[77] br[77] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_80 
+ bl[78] br[78] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_81 
+ bl[79] br[79] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_82 
+ bl[80] br[80] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_83 
+ bl[81] br[81] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_84 
+ bl[82] br[82] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_85 
+ bl[83] br[83] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_86 
+ bl[84] br[84] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_87 
+ bl[85] br[85] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_88 
+ bl[86] br[86] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_89 
+ bl[87] br[87] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_90 
+ bl[88] br[88] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_91 
+ bl[89] br[89] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_92 
+ bl[90] br[90] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_93 
+ bl[91] br[91] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_94 
+ bl[92] br[92] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_95 
+ bl[93] br[93] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_96 
+ bl[94] br[94] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_97 
+ bl[95] br[95] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_98 
+ bl[96] br[96] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_99 
+ bl[97] br[97] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_100 
+ bl[98] br[98] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_101 
+ bl[99] br[99] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_102 
+ bl[100] br[100] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_103 
+ bl[101] br[101] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_104 
+ bl[102] br[102] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_105 
+ bl[103] br[103] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_106 
+ bl[104] br[104] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_107 
+ bl[105] br[105] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_108 
+ bl[106] br[106] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_109 
+ bl[107] br[107] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_110 
+ bl[108] br[108] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_111 
+ bl[109] br[109] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_112 
+ bl[110] br[110] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_113 
+ bl[111] br[111] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_114 
+ bl[112] br[112] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_115 
+ bl[113] br[113] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_116 
+ bl[114] br[114] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_117 
+ bl[115] br[115] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_118 
+ bl[116] br[116] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_119 
+ bl[117] br[117] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_120 
+ bl[118] br[118] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_121 
+ bl[119] br[119] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_122 
+ bl[120] br[120] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_123 
+ bl[121] br[121] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_124 
+ bl[122] br[122] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_125 
+ bl[123] br[123] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_126 
+ bl[124] br[124] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_127 
+ bl[125] br[125] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_128 
+ bl[126] br[126] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_129 
+ bl[127] br[127] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_130 
+ vdd vdd vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_131 
+ vdd vdd vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_0 
+ vdd vdd vss vdd vpb vnb wl[12] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_14_1 
+ rbl rbr vss vdd vpb vnb wl[12] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_14_2 
+ bl[0] br[0] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_3 
+ bl[1] br[1] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_4 
+ bl[2] br[2] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_5 
+ bl[3] br[3] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_6 
+ bl[4] br[4] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_7 
+ bl[5] br[5] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_8 
+ bl[6] br[6] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_9 
+ bl[7] br[7] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_10 
+ bl[8] br[8] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_11 
+ bl[9] br[9] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_12 
+ bl[10] br[10] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_13 
+ bl[11] br[11] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_14 
+ bl[12] br[12] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_15 
+ bl[13] br[13] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_16 
+ bl[14] br[14] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_17 
+ bl[15] br[15] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_18 
+ bl[16] br[16] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_19 
+ bl[17] br[17] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_20 
+ bl[18] br[18] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_21 
+ bl[19] br[19] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_22 
+ bl[20] br[20] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_23 
+ bl[21] br[21] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_24 
+ bl[22] br[22] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_25 
+ bl[23] br[23] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_26 
+ bl[24] br[24] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_27 
+ bl[25] br[25] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_28 
+ bl[26] br[26] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_29 
+ bl[27] br[27] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_30 
+ bl[28] br[28] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_31 
+ bl[29] br[29] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_32 
+ bl[30] br[30] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_33 
+ bl[31] br[31] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_34 
+ bl[32] br[32] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_35 
+ bl[33] br[33] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_36 
+ bl[34] br[34] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_37 
+ bl[35] br[35] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_38 
+ bl[36] br[36] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_39 
+ bl[37] br[37] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_40 
+ bl[38] br[38] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_41 
+ bl[39] br[39] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_42 
+ bl[40] br[40] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_43 
+ bl[41] br[41] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_44 
+ bl[42] br[42] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_45 
+ bl[43] br[43] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_46 
+ bl[44] br[44] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_47 
+ bl[45] br[45] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_48 
+ bl[46] br[46] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_49 
+ bl[47] br[47] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_50 
+ bl[48] br[48] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_51 
+ bl[49] br[49] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_52 
+ bl[50] br[50] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_53 
+ bl[51] br[51] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_54 
+ bl[52] br[52] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_55 
+ bl[53] br[53] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_56 
+ bl[54] br[54] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_57 
+ bl[55] br[55] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_58 
+ bl[56] br[56] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_59 
+ bl[57] br[57] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_60 
+ bl[58] br[58] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_61 
+ bl[59] br[59] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_62 
+ bl[60] br[60] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_63 
+ bl[61] br[61] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_64 
+ bl[62] br[62] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_65 
+ bl[63] br[63] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_66 
+ bl[64] br[64] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_67 
+ bl[65] br[65] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_68 
+ bl[66] br[66] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_69 
+ bl[67] br[67] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_70 
+ bl[68] br[68] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_71 
+ bl[69] br[69] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_72 
+ bl[70] br[70] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_73 
+ bl[71] br[71] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_74 
+ bl[72] br[72] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_75 
+ bl[73] br[73] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_76 
+ bl[74] br[74] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_77 
+ bl[75] br[75] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_78 
+ bl[76] br[76] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_79 
+ bl[77] br[77] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_80 
+ bl[78] br[78] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_81 
+ bl[79] br[79] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_82 
+ bl[80] br[80] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_83 
+ bl[81] br[81] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_84 
+ bl[82] br[82] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_85 
+ bl[83] br[83] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_86 
+ bl[84] br[84] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_87 
+ bl[85] br[85] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_88 
+ bl[86] br[86] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_89 
+ bl[87] br[87] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_90 
+ bl[88] br[88] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_91 
+ bl[89] br[89] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_92 
+ bl[90] br[90] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_93 
+ bl[91] br[91] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_94 
+ bl[92] br[92] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_95 
+ bl[93] br[93] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_96 
+ bl[94] br[94] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_97 
+ bl[95] br[95] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_98 
+ bl[96] br[96] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_99 
+ bl[97] br[97] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_100 
+ bl[98] br[98] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_101 
+ bl[99] br[99] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_102 
+ bl[100] br[100] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_103 
+ bl[101] br[101] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_104 
+ bl[102] br[102] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_105 
+ bl[103] br[103] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_106 
+ bl[104] br[104] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_107 
+ bl[105] br[105] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_108 
+ bl[106] br[106] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_109 
+ bl[107] br[107] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_110 
+ bl[108] br[108] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_111 
+ bl[109] br[109] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_112 
+ bl[110] br[110] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_113 
+ bl[111] br[111] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_114 
+ bl[112] br[112] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_115 
+ bl[113] br[113] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_116 
+ bl[114] br[114] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_117 
+ bl[115] br[115] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_118 
+ bl[116] br[116] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_119 
+ bl[117] br[117] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_120 
+ bl[118] br[118] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_121 
+ bl[119] br[119] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_122 
+ bl[120] br[120] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_123 
+ bl[121] br[121] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_124 
+ bl[122] br[122] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_125 
+ bl[123] br[123] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_126 
+ bl[124] br[124] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_127 
+ bl[125] br[125] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_128 
+ bl[126] br[126] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_129 
+ bl[127] br[127] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_130 
+ vdd vdd vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_131 
+ vdd vdd vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_0 
+ vdd vdd vss vdd vpb vnb wl[13] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_15_1 
+ rbl rbr vss vdd vpb vnb wl[13] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_15_2 
+ bl[0] br[0] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_3 
+ bl[1] br[1] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_4 
+ bl[2] br[2] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_5 
+ bl[3] br[3] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_6 
+ bl[4] br[4] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_7 
+ bl[5] br[5] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_8 
+ bl[6] br[6] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_9 
+ bl[7] br[7] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_10 
+ bl[8] br[8] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_11 
+ bl[9] br[9] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_12 
+ bl[10] br[10] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_13 
+ bl[11] br[11] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_14 
+ bl[12] br[12] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_15 
+ bl[13] br[13] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_16 
+ bl[14] br[14] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_17 
+ bl[15] br[15] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_18 
+ bl[16] br[16] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_19 
+ bl[17] br[17] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_20 
+ bl[18] br[18] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_21 
+ bl[19] br[19] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_22 
+ bl[20] br[20] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_23 
+ bl[21] br[21] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_24 
+ bl[22] br[22] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_25 
+ bl[23] br[23] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_26 
+ bl[24] br[24] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_27 
+ bl[25] br[25] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_28 
+ bl[26] br[26] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_29 
+ bl[27] br[27] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_30 
+ bl[28] br[28] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_31 
+ bl[29] br[29] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_32 
+ bl[30] br[30] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_33 
+ bl[31] br[31] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_34 
+ bl[32] br[32] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_35 
+ bl[33] br[33] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_36 
+ bl[34] br[34] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_37 
+ bl[35] br[35] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_38 
+ bl[36] br[36] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_39 
+ bl[37] br[37] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_40 
+ bl[38] br[38] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_41 
+ bl[39] br[39] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_42 
+ bl[40] br[40] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_43 
+ bl[41] br[41] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_44 
+ bl[42] br[42] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_45 
+ bl[43] br[43] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_46 
+ bl[44] br[44] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_47 
+ bl[45] br[45] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_48 
+ bl[46] br[46] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_49 
+ bl[47] br[47] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_50 
+ bl[48] br[48] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_51 
+ bl[49] br[49] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_52 
+ bl[50] br[50] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_53 
+ bl[51] br[51] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_54 
+ bl[52] br[52] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_55 
+ bl[53] br[53] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_56 
+ bl[54] br[54] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_57 
+ bl[55] br[55] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_58 
+ bl[56] br[56] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_59 
+ bl[57] br[57] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_60 
+ bl[58] br[58] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_61 
+ bl[59] br[59] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_62 
+ bl[60] br[60] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_63 
+ bl[61] br[61] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_64 
+ bl[62] br[62] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_65 
+ bl[63] br[63] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_66 
+ bl[64] br[64] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_67 
+ bl[65] br[65] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_68 
+ bl[66] br[66] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_69 
+ bl[67] br[67] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_70 
+ bl[68] br[68] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_71 
+ bl[69] br[69] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_72 
+ bl[70] br[70] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_73 
+ bl[71] br[71] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_74 
+ bl[72] br[72] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_75 
+ bl[73] br[73] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_76 
+ bl[74] br[74] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_77 
+ bl[75] br[75] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_78 
+ bl[76] br[76] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_79 
+ bl[77] br[77] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_80 
+ bl[78] br[78] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_81 
+ bl[79] br[79] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_82 
+ bl[80] br[80] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_83 
+ bl[81] br[81] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_84 
+ bl[82] br[82] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_85 
+ bl[83] br[83] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_86 
+ bl[84] br[84] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_87 
+ bl[85] br[85] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_88 
+ bl[86] br[86] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_89 
+ bl[87] br[87] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_90 
+ bl[88] br[88] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_91 
+ bl[89] br[89] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_92 
+ bl[90] br[90] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_93 
+ bl[91] br[91] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_94 
+ bl[92] br[92] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_95 
+ bl[93] br[93] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_96 
+ bl[94] br[94] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_97 
+ bl[95] br[95] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_98 
+ bl[96] br[96] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_99 
+ bl[97] br[97] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_100 
+ bl[98] br[98] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_101 
+ bl[99] br[99] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_102 
+ bl[100] br[100] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_103 
+ bl[101] br[101] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_104 
+ bl[102] br[102] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_105 
+ bl[103] br[103] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_106 
+ bl[104] br[104] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_107 
+ bl[105] br[105] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_108 
+ bl[106] br[106] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_109 
+ bl[107] br[107] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_110 
+ bl[108] br[108] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_111 
+ bl[109] br[109] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_112 
+ bl[110] br[110] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_113 
+ bl[111] br[111] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_114 
+ bl[112] br[112] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_115 
+ bl[113] br[113] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_116 
+ bl[114] br[114] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_117 
+ bl[115] br[115] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_118 
+ bl[116] br[116] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_119 
+ bl[117] br[117] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_120 
+ bl[118] br[118] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_121 
+ bl[119] br[119] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_122 
+ bl[120] br[120] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_123 
+ bl[121] br[121] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_124 
+ bl[122] br[122] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_125 
+ bl[123] br[123] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_126 
+ bl[124] br[124] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_127 
+ bl[125] br[125] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_128 
+ bl[126] br[126] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_129 
+ bl[127] br[127] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_130 
+ vdd vdd vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_131 
+ vdd vdd vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_0 
+ vdd vdd vss vdd vpb vnb wl[14] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_16_1 
+ rbl rbr vss vdd vpb vnb wl[14] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_16_2 
+ bl[0] br[0] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_3 
+ bl[1] br[1] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_4 
+ bl[2] br[2] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_5 
+ bl[3] br[3] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_6 
+ bl[4] br[4] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_7 
+ bl[5] br[5] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_8 
+ bl[6] br[6] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_9 
+ bl[7] br[7] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_10 
+ bl[8] br[8] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_11 
+ bl[9] br[9] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_12 
+ bl[10] br[10] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_13 
+ bl[11] br[11] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_14 
+ bl[12] br[12] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_15 
+ bl[13] br[13] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_16 
+ bl[14] br[14] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_17 
+ bl[15] br[15] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_18 
+ bl[16] br[16] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_19 
+ bl[17] br[17] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_20 
+ bl[18] br[18] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_21 
+ bl[19] br[19] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_22 
+ bl[20] br[20] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_23 
+ bl[21] br[21] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_24 
+ bl[22] br[22] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_25 
+ bl[23] br[23] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_26 
+ bl[24] br[24] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_27 
+ bl[25] br[25] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_28 
+ bl[26] br[26] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_29 
+ bl[27] br[27] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_30 
+ bl[28] br[28] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_31 
+ bl[29] br[29] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_32 
+ bl[30] br[30] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_33 
+ bl[31] br[31] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_34 
+ bl[32] br[32] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_35 
+ bl[33] br[33] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_36 
+ bl[34] br[34] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_37 
+ bl[35] br[35] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_38 
+ bl[36] br[36] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_39 
+ bl[37] br[37] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_40 
+ bl[38] br[38] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_41 
+ bl[39] br[39] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_42 
+ bl[40] br[40] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_43 
+ bl[41] br[41] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_44 
+ bl[42] br[42] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_45 
+ bl[43] br[43] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_46 
+ bl[44] br[44] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_47 
+ bl[45] br[45] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_48 
+ bl[46] br[46] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_49 
+ bl[47] br[47] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_50 
+ bl[48] br[48] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_51 
+ bl[49] br[49] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_52 
+ bl[50] br[50] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_53 
+ bl[51] br[51] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_54 
+ bl[52] br[52] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_55 
+ bl[53] br[53] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_56 
+ bl[54] br[54] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_57 
+ bl[55] br[55] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_58 
+ bl[56] br[56] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_59 
+ bl[57] br[57] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_60 
+ bl[58] br[58] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_61 
+ bl[59] br[59] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_62 
+ bl[60] br[60] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_63 
+ bl[61] br[61] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_64 
+ bl[62] br[62] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_65 
+ bl[63] br[63] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_66 
+ bl[64] br[64] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_67 
+ bl[65] br[65] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_68 
+ bl[66] br[66] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_69 
+ bl[67] br[67] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_70 
+ bl[68] br[68] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_71 
+ bl[69] br[69] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_72 
+ bl[70] br[70] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_73 
+ bl[71] br[71] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_74 
+ bl[72] br[72] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_75 
+ bl[73] br[73] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_76 
+ bl[74] br[74] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_77 
+ bl[75] br[75] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_78 
+ bl[76] br[76] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_79 
+ bl[77] br[77] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_80 
+ bl[78] br[78] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_81 
+ bl[79] br[79] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_82 
+ bl[80] br[80] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_83 
+ bl[81] br[81] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_84 
+ bl[82] br[82] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_85 
+ bl[83] br[83] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_86 
+ bl[84] br[84] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_87 
+ bl[85] br[85] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_88 
+ bl[86] br[86] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_89 
+ bl[87] br[87] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_90 
+ bl[88] br[88] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_91 
+ bl[89] br[89] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_92 
+ bl[90] br[90] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_93 
+ bl[91] br[91] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_94 
+ bl[92] br[92] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_95 
+ bl[93] br[93] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_96 
+ bl[94] br[94] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_97 
+ bl[95] br[95] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_98 
+ bl[96] br[96] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_99 
+ bl[97] br[97] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_100 
+ bl[98] br[98] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_101 
+ bl[99] br[99] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_102 
+ bl[100] br[100] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_103 
+ bl[101] br[101] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_104 
+ bl[102] br[102] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_105 
+ bl[103] br[103] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_106 
+ bl[104] br[104] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_107 
+ bl[105] br[105] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_108 
+ bl[106] br[106] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_109 
+ bl[107] br[107] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_110 
+ bl[108] br[108] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_111 
+ bl[109] br[109] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_112 
+ bl[110] br[110] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_113 
+ bl[111] br[111] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_114 
+ bl[112] br[112] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_115 
+ bl[113] br[113] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_116 
+ bl[114] br[114] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_117 
+ bl[115] br[115] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_118 
+ bl[116] br[116] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_119 
+ bl[117] br[117] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_120 
+ bl[118] br[118] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_121 
+ bl[119] br[119] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_122 
+ bl[120] br[120] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_123 
+ bl[121] br[121] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_124 
+ bl[122] br[122] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_125 
+ bl[123] br[123] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_126 
+ bl[124] br[124] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_127 
+ bl[125] br[125] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_128 
+ bl[126] br[126] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_129 
+ bl[127] br[127] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_130 
+ vdd vdd vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_131 
+ vdd vdd vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_0 
+ vdd vdd vss vdd vpb vnb wl[15] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_17_1 
+ rbl rbr vss vdd vpb vnb wl[15] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_17_2 
+ bl[0] br[0] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_3 
+ bl[1] br[1] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_4 
+ bl[2] br[2] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_5 
+ bl[3] br[3] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_6 
+ bl[4] br[4] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_7 
+ bl[5] br[5] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_8 
+ bl[6] br[6] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_9 
+ bl[7] br[7] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_10 
+ bl[8] br[8] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_11 
+ bl[9] br[9] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_12 
+ bl[10] br[10] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_13 
+ bl[11] br[11] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_14 
+ bl[12] br[12] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_15 
+ bl[13] br[13] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_16 
+ bl[14] br[14] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_17 
+ bl[15] br[15] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_18 
+ bl[16] br[16] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_19 
+ bl[17] br[17] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_20 
+ bl[18] br[18] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_21 
+ bl[19] br[19] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_22 
+ bl[20] br[20] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_23 
+ bl[21] br[21] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_24 
+ bl[22] br[22] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_25 
+ bl[23] br[23] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_26 
+ bl[24] br[24] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_27 
+ bl[25] br[25] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_28 
+ bl[26] br[26] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_29 
+ bl[27] br[27] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_30 
+ bl[28] br[28] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_31 
+ bl[29] br[29] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_32 
+ bl[30] br[30] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_33 
+ bl[31] br[31] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_34 
+ bl[32] br[32] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_35 
+ bl[33] br[33] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_36 
+ bl[34] br[34] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_37 
+ bl[35] br[35] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_38 
+ bl[36] br[36] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_39 
+ bl[37] br[37] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_40 
+ bl[38] br[38] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_41 
+ bl[39] br[39] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_42 
+ bl[40] br[40] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_43 
+ bl[41] br[41] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_44 
+ bl[42] br[42] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_45 
+ bl[43] br[43] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_46 
+ bl[44] br[44] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_47 
+ bl[45] br[45] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_48 
+ bl[46] br[46] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_49 
+ bl[47] br[47] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_50 
+ bl[48] br[48] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_51 
+ bl[49] br[49] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_52 
+ bl[50] br[50] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_53 
+ bl[51] br[51] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_54 
+ bl[52] br[52] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_55 
+ bl[53] br[53] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_56 
+ bl[54] br[54] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_57 
+ bl[55] br[55] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_58 
+ bl[56] br[56] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_59 
+ bl[57] br[57] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_60 
+ bl[58] br[58] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_61 
+ bl[59] br[59] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_62 
+ bl[60] br[60] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_63 
+ bl[61] br[61] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_64 
+ bl[62] br[62] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_65 
+ bl[63] br[63] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_66 
+ bl[64] br[64] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_67 
+ bl[65] br[65] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_68 
+ bl[66] br[66] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_69 
+ bl[67] br[67] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_70 
+ bl[68] br[68] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_71 
+ bl[69] br[69] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_72 
+ bl[70] br[70] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_73 
+ bl[71] br[71] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_74 
+ bl[72] br[72] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_75 
+ bl[73] br[73] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_76 
+ bl[74] br[74] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_77 
+ bl[75] br[75] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_78 
+ bl[76] br[76] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_79 
+ bl[77] br[77] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_80 
+ bl[78] br[78] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_81 
+ bl[79] br[79] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_82 
+ bl[80] br[80] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_83 
+ bl[81] br[81] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_84 
+ bl[82] br[82] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_85 
+ bl[83] br[83] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_86 
+ bl[84] br[84] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_87 
+ bl[85] br[85] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_88 
+ bl[86] br[86] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_89 
+ bl[87] br[87] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_90 
+ bl[88] br[88] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_91 
+ bl[89] br[89] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_92 
+ bl[90] br[90] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_93 
+ bl[91] br[91] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_94 
+ bl[92] br[92] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_95 
+ bl[93] br[93] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_96 
+ bl[94] br[94] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_97 
+ bl[95] br[95] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_98 
+ bl[96] br[96] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_99 
+ bl[97] br[97] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_100 
+ bl[98] br[98] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_101 
+ bl[99] br[99] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_102 
+ bl[100] br[100] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_103 
+ bl[101] br[101] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_104 
+ bl[102] br[102] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_105 
+ bl[103] br[103] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_106 
+ bl[104] br[104] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_107 
+ bl[105] br[105] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_108 
+ bl[106] br[106] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_109 
+ bl[107] br[107] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_110 
+ bl[108] br[108] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_111 
+ bl[109] br[109] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_112 
+ bl[110] br[110] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_113 
+ bl[111] br[111] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_114 
+ bl[112] br[112] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_115 
+ bl[113] br[113] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_116 
+ bl[114] br[114] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_117 
+ bl[115] br[115] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_118 
+ bl[116] br[116] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_119 
+ bl[117] br[117] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_120 
+ bl[118] br[118] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_121 
+ bl[119] br[119] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_122 
+ bl[120] br[120] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_123 
+ bl[121] br[121] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_124 
+ bl[122] br[122] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_125 
+ bl[123] br[123] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_126 
+ bl[124] br[124] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_127 
+ bl[125] br[125] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_128 
+ bl[126] br[126] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_129 
+ bl[127] br[127] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_130 
+ vdd vdd vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_131 
+ vdd vdd vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_0 
+ vdd vdd vss vdd vpb vnb wl[16] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_18_1 
+ rbl rbr vss vdd vpb vnb wl[16] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_18_2 
+ bl[0] br[0] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_3 
+ bl[1] br[1] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_4 
+ bl[2] br[2] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_5 
+ bl[3] br[3] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_6 
+ bl[4] br[4] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_7 
+ bl[5] br[5] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_8 
+ bl[6] br[6] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_9 
+ bl[7] br[7] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_10 
+ bl[8] br[8] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_11 
+ bl[9] br[9] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_12 
+ bl[10] br[10] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_13 
+ bl[11] br[11] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_14 
+ bl[12] br[12] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_15 
+ bl[13] br[13] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_16 
+ bl[14] br[14] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_17 
+ bl[15] br[15] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_18 
+ bl[16] br[16] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_19 
+ bl[17] br[17] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_20 
+ bl[18] br[18] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_21 
+ bl[19] br[19] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_22 
+ bl[20] br[20] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_23 
+ bl[21] br[21] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_24 
+ bl[22] br[22] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_25 
+ bl[23] br[23] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_26 
+ bl[24] br[24] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_27 
+ bl[25] br[25] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_28 
+ bl[26] br[26] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_29 
+ bl[27] br[27] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_30 
+ bl[28] br[28] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_31 
+ bl[29] br[29] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_32 
+ bl[30] br[30] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_33 
+ bl[31] br[31] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_34 
+ bl[32] br[32] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_35 
+ bl[33] br[33] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_36 
+ bl[34] br[34] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_37 
+ bl[35] br[35] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_38 
+ bl[36] br[36] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_39 
+ bl[37] br[37] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_40 
+ bl[38] br[38] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_41 
+ bl[39] br[39] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_42 
+ bl[40] br[40] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_43 
+ bl[41] br[41] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_44 
+ bl[42] br[42] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_45 
+ bl[43] br[43] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_46 
+ bl[44] br[44] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_47 
+ bl[45] br[45] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_48 
+ bl[46] br[46] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_49 
+ bl[47] br[47] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_50 
+ bl[48] br[48] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_51 
+ bl[49] br[49] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_52 
+ bl[50] br[50] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_53 
+ bl[51] br[51] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_54 
+ bl[52] br[52] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_55 
+ bl[53] br[53] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_56 
+ bl[54] br[54] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_57 
+ bl[55] br[55] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_58 
+ bl[56] br[56] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_59 
+ bl[57] br[57] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_60 
+ bl[58] br[58] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_61 
+ bl[59] br[59] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_62 
+ bl[60] br[60] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_63 
+ bl[61] br[61] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_64 
+ bl[62] br[62] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_65 
+ bl[63] br[63] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_66 
+ bl[64] br[64] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_67 
+ bl[65] br[65] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_68 
+ bl[66] br[66] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_69 
+ bl[67] br[67] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_70 
+ bl[68] br[68] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_71 
+ bl[69] br[69] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_72 
+ bl[70] br[70] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_73 
+ bl[71] br[71] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_74 
+ bl[72] br[72] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_75 
+ bl[73] br[73] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_76 
+ bl[74] br[74] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_77 
+ bl[75] br[75] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_78 
+ bl[76] br[76] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_79 
+ bl[77] br[77] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_80 
+ bl[78] br[78] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_81 
+ bl[79] br[79] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_82 
+ bl[80] br[80] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_83 
+ bl[81] br[81] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_84 
+ bl[82] br[82] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_85 
+ bl[83] br[83] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_86 
+ bl[84] br[84] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_87 
+ bl[85] br[85] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_88 
+ bl[86] br[86] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_89 
+ bl[87] br[87] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_90 
+ bl[88] br[88] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_91 
+ bl[89] br[89] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_92 
+ bl[90] br[90] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_93 
+ bl[91] br[91] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_94 
+ bl[92] br[92] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_95 
+ bl[93] br[93] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_96 
+ bl[94] br[94] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_97 
+ bl[95] br[95] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_98 
+ bl[96] br[96] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_99 
+ bl[97] br[97] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_100 
+ bl[98] br[98] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_101 
+ bl[99] br[99] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_102 
+ bl[100] br[100] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_103 
+ bl[101] br[101] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_104 
+ bl[102] br[102] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_105 
+ bl[103] br[103] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_106 
+ bl[104] br[104] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_107 
+ bl[105] br[105] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_108 
+ bl[106] br[106] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_109 
+ bl[107] br[107] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_110 
+ bl[108] br[108] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_111 
+ bl[109] br[109] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_112 
+ bl[110] br[110] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_113 
+ bl[111] br[111] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_114 
+ bl[112] br[112] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_115 
+ bl[113] br[113] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_116 
+ bl[114] br[114] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_117 
+ bl[115] br[115] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_118 
+ bl[116] br[116] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_119 
+ bl[117] br[117] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_120 
+ bl[118] br[118] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_121 
+ bl[119] br[119] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_122 
+ bl[120] br[120] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_123 
+ bl[121] br[121] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_124 
+ bl[122] br[122] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_125 
+ bl[123] br[123] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_126 
+ bl[124] br[124] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_127 
+ bl[125] br[125] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_128 
+ bl[126] br[126] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_129 
+ bl[127] br[127] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_130 
+ vdd vdd vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_131 
+ vdd vdd vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_0 
+ vdd vdd vss vdd vpb vnb wl[17] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_19_1 
+ rbl rbr vss vdd vpb vnb wl[17] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_19_2 
+ bl[0] br[0] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_3 
+ bl[1] br[1] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_4 
+ bl[2] br[2] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_5 
+ bl[3] br[3] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_6 
+ bl[4] br[4] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_7 
+ bl[5] br[5] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_8 
+ bl[6] br[6] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_9 
+ bl[7] br[7] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_10 
+ bl[8] br[8] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_11 
+ bl[9] br[9] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_12 
+ bl[10] br[10] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_13 
+ bl[11] br[11] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_14 
+ bl[12] br[12] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_15 
+ bl[13] br[13] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_16 
+ bl[14] br[14] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_17 
+ bl[15] br[15] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_18 
+ bl[16] br[16] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_19 
+ bl[17] br[17] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_20 
+ bl[18] br[18] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_21 
+ bl[19] br[19] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_22 
+ bl[20] br[20] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_23 
+ bl[21] br[21] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_24 
+ bl[22] br[22] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_25 
+ bl[23] br[23] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_26 
+ bl[24] br[24] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_27 
+ bl[25] br[25] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_28 
+ bl[26] br[26] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_29 
+ bl[27] br[27] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_30 
+ bl[28] br[28] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_31 
+ bl[29] br[29] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_32 
+ bl[30] br[30] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_33 
+ bl[31] br[31] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_34 
+ bl[32] br[32] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_35 
+ bl[33] br[33] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_36 
+ bl[34] br[34] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_37 
+ bl[35] br[35] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_38 
+ bl[36] br[36] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_39 
+ bl[37] br[37] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_40 
+ bl[38] br[38] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_41 
+ bl[39] br[39] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_42 
+ bl[40] br[40] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_43 
+ bl[41] br[41] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_44 
+ bl[42] br[42] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_45 
+ bl[43] br[43] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_46 
+ bl[44] br[44] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_47 
+ bl[45] br[45] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_48 
+ bl[46] br[46] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_49 
+ bl[47] br[47] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_50 
+ bl[48] br[48] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_51 
+ bl[49] br[49] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_52 
+ bl[50] br[50] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_53 
+ bl[51] br[51] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_54 
+ bl[52] br[52] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_55 
+ bl[53] br[53] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_56 
+ bl[54] br[54] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_57 
+ bl[55] br[55] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_58 
+ bl[56] br[56] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_59 
+ bl[57] br[57] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_60 
+ bl[58] br[58] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_61 
+ bl[59] br[59] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_62 
+ bl[60] br[60] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_63 
+ bl[61] br[61] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_64 
+ bl[62] br[62] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_65 
+ bl[63] br[63] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_66 
+ bl[64] br[64] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_67 
+ bl[65] br[65] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_68 
+ bl[66] br[66] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_69 
+ bl[67] br[67] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_70 
+ bl[68] br[68] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_71 
+ bl[69] br[69] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_72 
+ bl[70] br[70] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_73 
+ bl[71] br[71] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_74 
+ bl[72] br[72] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_75 
+ bl[73] br[73] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_76 
+ bl[74] br[74] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_77 
+ bl[75] br[75] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_78 
+ bl[76] br[76] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_79 
+ bl[77] br[77] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_80 
+ bl[78] br[78] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_81 
+ bl[79] br[79] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_82 
+ bl[80] br[80] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_83 
+ bl[81] br[81] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_84 
+ bl[82] br[82] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_85 
+ bl[83] br[83] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_86 
+ bl[84] br[84] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_87 
+ bl[85] br[85] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_88 
+ bl[86] br[86] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_89 
+ bl[87] br[87] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_90 
+ bl[88] br[88] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_91 
+ bl[89] br[89] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_92 
+ bl[90] br[90] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_93 
+ bl[91] br[91] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_94 
+ bl[92] br[92] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_95 
+ bl[93] br[93] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_96 
+ bl[94] br[94] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_97 
+ bl[95] br[95] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_98 
+ bl[96] br[96] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_99 
+ bl[97] br[97] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_100 
+ bl[98] br[98] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_101 
+ bl[99] br[99] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_102 
+ bl[100] br[100] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_103 
+ bl[101] br[101] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_104 
+ bl[102] br[102] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_105 
+ bl[103] br[103] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_106 
+ bl[104] br[104] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_107 
+ bl[105] br[105] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_108 
+ bl[106] br[106] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_109 
+ bl[107] br[107] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_110 
+ bl[108] br[108] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_111 
+ bl[109] br[109] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_112 
+ bl[110] br[110] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_113 
+ bl[111] br[111] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_114 
+ bl[112] br[112] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_115 
+ bl[113] br[113] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_116 
+ bl[114] br[114] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_117 
+ bl[115] br[115] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_118 
+ bl[116] br[116] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_119 
+ bl[117] br[117] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_120 
+ bl[118] br[118] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_121 
+ bl[119] br[119] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_122 
+ bl[120] br[120] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_123 
+ bl[121] br[121] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_124 
+ bl[122] br[122] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_125 
+ bl[123] br[123] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_126 
+ bl[124] br[124] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_127 
+ bl[125] br[125] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_128 
+ bl[126] br[126] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_129 
+ bl[127] br[127] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_130 
+ vdd vdd vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_131 
+ vdd vdd vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_0 
+ vdd vdd vss vdd vpb vnb wl[18] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_20_1 
+ rbl rbr vss vdd vpb vnb wl[18] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_20_2 
+ bl[0] br[0] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_3 
+ bl[1] br[1] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_4 
+ bl[2] br[2] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_5 
+ bl[3] br[3] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_6 
+ bl[4] br[4] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_7 
+ bl[5] br[5] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_8 
+ bl[6] br[6] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_9 
+ bl[7] br[7] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_10 
+ bl[8] br[8] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_11 
+ bl[9] br[9] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_12 
+ bl[10] br[10] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_13 
+ bl[11] br[11] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_14 
+ bl[12] br[12] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_15 
+ bl[13] br[13] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_16 
+ bl[14] br[14] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_17 
+ bl[15] br[15] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_18 
+ bl[16] br[16] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_19 
+ bl[17] br[17] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_20 
+ bl[18] br[18] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_21 
+ bl[19] br[19] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_22 
+ bl[20] br[20] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_23 
+ bl[21] br[21] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_24 
+ bl[22] br[22] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_25 
+ bl[23] br[23] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_26 
+ bl[24] br[24] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_27 
+ bl[25] br[25] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_28 
+ bl[26] br[26] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_29 
+ bl[27] br[27] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_30 
+ bl[28] br[28] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_31 
+ bl[29] br[29] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_32 
+ bl[30] br[30] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_33 
+ bl[31] br[31] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_34 
+ bl[32] br[32] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_35 
+ bl[33] br[33] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_36 
+ bl[34] br[34] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_37 
+ bl[35] br[35] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_38 
+ bl[36] br[36] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_39 
+ bl[37] br[37] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_40 
+ bl[38] br[38] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_41 
+ bl[39] br[39] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_42 
+ bl[40] br[40] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_43 
+ bl[41] br[41] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_44 
+ bl[42] br[42] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_45 
+ bl[43] br[43] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_46 
+ bl[44] br[44] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_47 
+ bl[45] br[45] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_48 
+ bl[46] br[46] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_49 
+ bl[47] br[47] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_50 
+ bl[48] br[48] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_51 
+ bl[49] br[49] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_52 
+ bl[50] br[50] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_53 
+ bl[51] br[51] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_54 
+ bl[52] br[52] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_55 
+ bl[53] br[53] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_56 
+ bl[54] br[54] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_57 
+ bl[55] br[55] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_58 
+ bl[56] br[56] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_59 
+ bl[57] br[57] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_60 
+ bl[58] br[58] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_61 
+ bl[59] br[59] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_62 
+ bl[60] br[60] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_63 
+ bl[61] br[61] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_64 
+ bl[62] br[62] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_65 
+ bl[63] br[63] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_66 
+ bl[64] br[64] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_67 
+ bl[65] br[65] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_68 
+ bl[66] br[66] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_69 
+ bl[67] br[67] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_70 
+ bl[68] br[68] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_71 
+ bl[69] br[69] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_72 
+ bl[70] br[70] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_73 
+ bl[71] br[71] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_74 
+ bl[72] br[72] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_75 
+ bl[73] br[73] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_76 
+ bl[74] br[74] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_77 
+ bl[75] br[75] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_78 
+ bl[76] br[76] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_79 
+ bl[77] br[77] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_80 
+ bl[78] br[78] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_81 
+ bl[79] br[79] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_82 
+ bl[80] br[80] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_83 
+ bl[81] br[81] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_84 
+ bl[82] br[82] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_85 
+ bl[83] br[83] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_86 
+ bl[84] br[84] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_87 
+ bl[85] br[85] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_88 
+ bl[86] br[86] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_89 
+ bl[87] br[87] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_90 
+ bl[88] br[88] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_91 
+ bl[89] br[89] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_92 
+ bl[90] br[90] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_93 
+ bl[91] br[91] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_94 
+ bl[92] br[92] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_95 
+ bl[93] br[93] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_96 
+ bl[94] br[94] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_97 
+ bl[95] br[95] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_98 
+ bl[96] br[96] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_99 
+ bl[97] br[97] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_100 
+ bl[98] br[98] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_101 
+ bl[99] br[99] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_102 
+ bl[100] br[100] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_103 
+ bl[101] br[101] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_104 
+ bl[102] br[102] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_105 
+ bl[103] br[103] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_106 
+ bl[104] br[104] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_107 
+ bl[105] br[105] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_108 
+ bl[106] br[106] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_109 
+ bl[107] br[107] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_110 
+ bl[108] br[108] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_111 
+ bl[109] br[109] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_112 
+ bl[110] br[110] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_113 
+ bl[111] br[111] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_114 
+ bl[112] br[112] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_115 
+ bl[113] br[113] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_116 
+ bl[114] br[114] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_117 
+ bl[115] br[115] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_118 
+ bl[116] br[116] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_119 
+ bl[117] br[117] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_120 
+ bl[118] br[118] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_121 
+ bl[119] br[119] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_122 
+ bl[120] br[120] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_123 
+ bl[121] br[121] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_124 
+ bl[122] br[122] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_125 
+ bl[123] br[123] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_126 
+ bl[124] br[124] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_127 
+ bl[125] br[125] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_128 
+ bl[126] br[126] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_129 
+ bl[127] br[127] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_130 
+ vdd vdd vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_131 
+ vdd vdd vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_0 
+ vdd vdd vss vdd vpb vnb wl[19] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_21_1 
+ rbl rbr vss vdd vpb vnb wl[19] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_21_2 
+ bl[0] br[0] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_3 
+ bl[1] br[1] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_4 
+ bl[2] br[2] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_5 
+ bl[3] br[3] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_6 
+ bl[4] br[4] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_7 
+ bl[5] br[5] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_8 
+ bl[6] br[6] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_9 
+ bl[7] br[7] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_10 
+ bl[8] br[8] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_11 
+ bl[9] br[9] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_12 
+ bl[10] br[10] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_13 
+ bl[11] br[11] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_14 
+ bl[12] br[12] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_15 
+ bl[13] br[13] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_16 
+ bl[14] br[14] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_17 
+ bl[15] br[15] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_18 
+ bl[16] br[16] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_19 
+ bl[17] br[17] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_20 
+ bl[18] br[18] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_21 
+ bl[19] br[19] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_22 
+ bl[20] br[20] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_23 
+ bl[21] br[21] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_24 
+ bl[22] br[22] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_25 
+ bl[23] br[23] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_26 
+ bl[24] br[24] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_27 
+ bl[25] br[25] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_28 
+ bl[26] br[26] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_29 
+ bl[27] br[27] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_30 
+ bl[28] br[28] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_31 
+ bl[29] br[29] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_32 
+ bl[30] br[30] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_33 
+ bl[31] br[31] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_34 
+ bl[32] br[32] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_35 
+ bl[33] br[33] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_36 
+ bl[34] br[34] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_37 
+ bl[35] br[35] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_38 
+ bl[36] br[36] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_39 
+ bl[37] br[37] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_40 
+ bl[38] br[38] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_41 
+ bl[39] br[39] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_42 
+ bl[40] br[40] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_43 
+ bl[41] br[41] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_44 
+ bl[42] br[42] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_45 
+ bl[43] br[43] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_46 
+ bl[44] br[44] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_47 
+ bl[45] br[45] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_48 
+ bl[46] br[46] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_49 
+ bl[47] br[47] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_50 
+ bl[48] br[48] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_51 
+ bl[49] br[49] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_52 
+ bl[50] br[50] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_53 
+ bl[51] br[51] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_54 
+ bl[52] br[52] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_55 
+ bl[53] br[53] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_56 
+ bl[54] br[54] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_57 
+ bl[55] br[55] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_58 
+ bl[56] br[56] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_59 
+ bl[57] br[57] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_60 
+ bl[58] br[58] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_61 
+ bl[59] br[59] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_62 
+ bl[60] br[60] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_63 
+ bl[61] br[61] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_64 
+ bl[62] br[62] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_65 
+ bl[63] br[63] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_66 
+ bl[64] br[64] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_67 
+ bl[65] br[65] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_68 
+ bl[66] br[66] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_69 
+ bl[67] br[67] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_70 
+ bl[68] br[68] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_71 
+ bl[69] br[69] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_72 
+ bl[70] br[70] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_73 
+ bl[71] br[71] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_74 
+ bl[72] br[72] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_75 
+ bl[73] br[73] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_76 
+ bl[74] br[74] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_77 
+ bl[75] br[75] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_78 
+ bl[76] br[76] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_79 
+ bl[77] br[77] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_80 
+ bl[78] br[78] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_81 
+ bl[79] br[79] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_82 
+ bl[80] br[80] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_83 
+ bl[81] br[81] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_84 
+ bl[82] br[82] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_85 
+ bl[83] br[83] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_86 
+ bl[84] br[84] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_87 
+ bl[85] br[85] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_88 
+ bl[86] br[86] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_89 
+ bl[87] br[87] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_90 
+ bl[88] br[88] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_91 
+ bl[89] br[89] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_92 
+ bl[90] br[90] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_93 
+ bl[91] br[91] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_94 
+ bl[92] br[92] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_95 
+ bl[93] br[93] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_96 
+ bl[94] br[94] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_97 
+ bl[95] br[95] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_98 
+ bl[96] br[96] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_99 
+ bl[97] br[97] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_100 
+ bl[98] br[98] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_101 
+ bl[99] br[99] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_102 
+ bl[100] br[100] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_103 
+ bl[101] br[101] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_104 
+ bl[102] br[102] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_105 
+ bl[103] br[103] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_106 
+ bl[104] br[104] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_107 
+ bl[105] br[105] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_108 
+ bl[106] br[106] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_109 
+ bl[107] br[107] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_110 
+ bl[108] br[108] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_111 
+ bl[109] br[109] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_112 
+ bl[110] br[110] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_113 
+ bl[111] br[111] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_114 
+ bl[112] br[112] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_115 
+ bl[113] br[113] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_116 
+ bl[114] br[114] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_117 
+ bl[115] br[115] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_118 
+ bl[116] br[116] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_119 
+ bl[117] br[117] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_120 
+ bl[118] br[118] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_121 
+ bl[119] br[119] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_122 
+ bl[120] br[120] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_123 
+ bl[121] br[121] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_124 
+ bl[122] br[122] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_125 
+ bl[123] br[123] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_126 
+ bl[124] br[124] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_127 
+ bl[125] br[125] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_128 
+ bl[126] br[126] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_129 
+ bl[127] br[127] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_130 
+ vdd vdd vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_131 
+ vdd vdd vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_0 
+ vdd vdd vss vdd vpb vnb wl[20] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_22_1 
+ rbl rbr vss vdd vpb vnb wl[20] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_22_2 
+ bl[0] br[0] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_3 
+ bl[1] br[1] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_4 
+ bl[2] br[2] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_5 
+ bl[3] br[3] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_6 
+ bl[4] br[4] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_7 
+ bl[5] br[5] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_8 
+ bl[6] br[6] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_9 
+ bl[7] br[7] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_10 
+ bl[8] br[8] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_11 
+ bl[9] br[9] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_12 
+ bl[10] br[10] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_13 
+ bl[11] br[11] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_14 
+ bl[12] br[12] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_15 
+ bl[13] br[13] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_16 
+ bl[14] br[14] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_17 
+ bl[15] br[15] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_18 
+ bl[16] br[16] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_19 
+ bl[17] br[17] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_20 
+ bl[18] br[18] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_21 
+ bl[19] br[19] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_22 
+ bl[20] br[20] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_23 
+ bl[21] br[21] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_24 
+ bl[22] br[22] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_25 
+ bl[23] br[23] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_26 
+ bl[24] br[24] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_27 
+ bl[25] br[25] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_28 
+ bl[26] br[26] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_29 
+ bl[27] br[27] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_30 
+ bl[28] br[28] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_31 
+ bl[29] br[29] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_32 
+ bl[30] br[30] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_33 
+ bl[31] br[31] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_34 
+ bl[32] br[32] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_35 
+ bl[33] br[33] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_36 
+ bl[34] br[34] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_37 
+ bl[35] br[35] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_38 
+ bl[36] br[36] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_39 
+ bl[37] br[37] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_40 
+ bl[38] br[38] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_41 
+ bl[39] br[39] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_42 
+ bl[40] br[40] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_43 
+ bl[41] br[41] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_44 
+ bl[42] br[42] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_45 
+ bl[43] br[43] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_46 
+ bl[44] br[44] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_47 
+ bl[45] br[45] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_48 
+ bl[46] br[46] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_49 
+ bl[47] br[47] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_50 
+ bl[48] br[48] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_51 
+ bl[49] br[49] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_52 
+ bl[50] br[50] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_53 
+ bl[51] br[51] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_54 
+ bl[52] br[52] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_55 
+ bl[53] br[53] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_56 
+ bl[54] br[54] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_57 
+ bl[55] br[55] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_58 
+ bl[56] br[56] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_59 
+ bl[57] br[57] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_60 
+ bl[58] br[58] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_61 
+ bl[59] br[59] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_62 
+ bl[60] br[60] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_63 
+ bl[61] br[61] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_64 
+ bl[62] br[62] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_65 
+ bl[63] br[63] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_66 
+ bl[64] br[64] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_67 
+ bl[65] br[65] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_68 
+ bl[66] br[66] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_69 
+ bl[67] br[67] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_70 
+ bl[68] br[68] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_71 
+ bl[69] br[69] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_72 
+ bl[70] br[70] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_73 
+ bl[71] br[71] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_74 
+ bl[72] br[72] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_75 
+ bl[73] br[73] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_76 
+ bl[74] br[74] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_77 
+ bl[75] br[75] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_78 
+ bl[76] br[76] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_79 
+ bl[77] br[77] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_80 
+ bl[78] br[78] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_81 
+ bl[79] br[79] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_82 
+ bl[80] br[80] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_83 
+ bl[81] br[81] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_84 
+ bl[82] br[82] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_85 
+ bl[83] br[83] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_86 
+ bl[84] br[84] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_87 
+ bl[85] br[85] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_88 
+ bl[86] br[86] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_89 
+ bl[87] br[87] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_90 
+ bl[88] br[88] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_91 
+ bl[89] br[89] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_92 
+ bl[90] br[90] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_93 
+ bl[91] br[91] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_94 
+ bl[92] br[92] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_95 
+ bl[93] br[93] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_96 
+ bl[94] br[94] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_97 
+ bl[95] br[95] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_98 
+ bl[96] br[96] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_99 
+ bl[97] br[97] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_100 
+ bl[98] br[98] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_101 
+ bl[99] br[99] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_102 
+ bl[100] br[100] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_103 
+ bl[101] br[101] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_104 
+ bl[102] br[102] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_105 
+ bl[103] br[103] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_106 
+ bl[104] br[104] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_107 
+ bl[105] br[105] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_108 
+ bl[106] br[106] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_109 
+ bl[107] br[107] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_110 
+ bl[108] br[108] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_111 
+ bl[109] br[109] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_112 
+ bl[110] br[110] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_113 
+ bl[111] br[111] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_114 
+ bl[112] br[112] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_115 
+ bl[113] br[113] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_116 
+ bl[114] br[114] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_117 
+ bl[115] br[115] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_118 
+ bl[116] br[116] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_119 
+ bl[117] br[117] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_120 
+ bl[118] br[118] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_121 
+ bl[119] br[119] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_122 
+ bl[120] br[120] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_123 
+ bl[121] br[121] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_124 
+ bl[122] br[122] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_125 
+ bl[123] br[123] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_126 
+ bl[124] br[124] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_127 
+ bl[125] br[125] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_128 
+ bl[126] br[126] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_129 
+ bl[127] br[127] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_130 
+ vdd vdd vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_131 
+ vdd vdd vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_0 
+ vdd vdd vss vdd vpb vnb wl[21] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_23_1 
+ rbl rbr vss vdd vpb vnb wl[21] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_23_2 
+ bl[0] br[0] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_3 
+ bl[1] br[1] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_4 
+ bl[2] br[2] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_5 
+ bl[3] br[3] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_6 
+ bl[4] br[4] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_7 
+ bl[5] br[5] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_8 
+ bl[6] br[6] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_9 
+ bl[7] br[7] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_10 
+ bl[8] br[8] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_11 
+ bl[9] br[9] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_12 
+ bl[10] br[10] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_13 
+ bl[11] br[11] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_14 
+ bl[12] br[12] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_15 
+ bl[13] br[13] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_16 
+ bl[14] br[14] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_17 
+ bl[15] br[15] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_18 
+ bl[16] br[16] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_19 
+ bl[17] br[17] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_20 
+ bl[18] br[18] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_21 
+ bl[19] br[19] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_22 
+ bl[20] br[20] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_23 
+ bl[21] br[21] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_24 
+ bl[22] br[22] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_25 
+ bl[23] br[23] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_26 
+ bl[24] br[24] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_27 
+ bl[25] br[25] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_28 
+ bl[26] br[26] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_29 
+ bl[27] br[27] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_30 
+ bl[28] br[28] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_31 
+ bl[29] br[29] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_32 
+ bl[30] br[30] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_33 
+ bl[31] br[31] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_34 
+ bl[32] br[32] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_35 
+ bl[33] br[33] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_36 
+ bl[34] br[34] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_37 
+ bl[35] br[35] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_38 
+ bl[36] br[36] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_39 
+ bl[37] br[37] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_40 
+ bl[38] br[38] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_41 
+ bl[39] br[39] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_42 
+ bl[40] br[40] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_43 
+ bl[41] br[41] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_44 
+ bl[42] br[42] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_45 
+ bl[43] br[43] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_46 
+ bl[44] br[44] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_47 
+ bl[45] br[45] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_48 
+ bl[46] br[46] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_49 
+ bl[47] br[47] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_50 
+ bl[48] br[48] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_51 
+ bl[49] br[49] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_52 
+ bl[50] br[50] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_53 
+ bl[51] br[51] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_54 
+ bl[52] br[52] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_55 
+ bl[53] br[53] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_56 
+ bl[54] br[54] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_57 
+ bl[55] br[55] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_58 
+ bl[56] br[56] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_59 
+ bl[57] br[57] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_60 
+ bl[58] br[58] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_61 
+ bl[59] br[59] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_62 
+ bl[60] br[60] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_63 
+ bl[61] br[61] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_64 
+ bl[62] br[62] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_65 
+ bl[63] br[63] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_66 
+ bl[64] br[64] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_67 
+ bl[65] br[65] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_68 
+ bl[66] br[66] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_69 
+ bl[67] br[67] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_70 
+ bl[68] br[68] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_71 
+ bl[69] br[69] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_72 
+ bl[70] br[70] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_73 
+ bl[71] br[71] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_74 
+ bl[72] br[72] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_75 
+ bl[73] br[73] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_76 
+ bl[74] br[74] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_77 
+ bl[75] br[75] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_78 
+ bl[76] br[76] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_79 
+ bl[77] br[77] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_80 
+ bl[78] br[78] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_81 
+ bl[79] br[79] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_82 
+ bl[80] br[80] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_83 
+ bl[81] br[81] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_84 
+ bl[82] br[82] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_85 
+ bl[83] br[83] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_86 
+ bl[84] br[84] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_87 
+ bl[85] br[85] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_88 
+ bl[86] br[86] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_89 
+ bl[87] br[87] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_90 
+ bl[88] br[88] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_91 
+ bl[89] br[89] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_92 
+ bl[90] br[90] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_93 
+ bl[91] br[91] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_94 
+ bl[92] br[92] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_95 
+ bl[93] br[93] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_96 
+ bl[94] br[94] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_97 
+ bl[95] br[95] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_98 
+ bl[96] br[96] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_99 
+ bl[97] br[97] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_100 
+ bl[98] br[98] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_101 
+ bl[99] br[99] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_102 
+ bl[100] br[100] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_103 
+ bl[101] br[101] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_104 
+ bl[102] br[102] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_105 
+ bl[103] br[103] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_106 
+ bl[104] br[104] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_107 
+ bl[105] br[105] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_108 
+ bl[106] br[106] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_109 
+ bl[107] br[107] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_110 
+ bl[108] br[108] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_111 
+ bl[109] br[109] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_112 
+ bl[110] br[110] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_113 
+ bl[111] br[111] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_114 
+ bl[112] br[112] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_115 
+ bl[113] br[113] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_116 
+ bl[114] br[114] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_117 
+ bl[115] br[115] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_118 
+ bl[116] br[116] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_119 
+ bl[117] br[117] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_120 
+ bl[118] br[118] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_121 
+ bl[119] br[119] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_122 
+ bl[120] br[120] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_123 
+ bl[121] br[121] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_124 
+ bl[122] br[122] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_125 
+ bl[123] br[123] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_126 
+ bl[124] br[124] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_127 
+ bl[125] br[125] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_128 
+ bl[126] br[126] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_129 
+ bl[127] br[127] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_130 
+ vdd vdd vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_131 
+ vdd vdd vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_0 
+ vdd vdd vss vdd vpb vnb wl[22] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_24_1 
+ rbl rbr vss vdd vpb vnb wl[22] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_24_2 
+ bl[0] br[0] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_3 
+ bl[1] br[1] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_4 
+ bl[2] br[2] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_5 
+ bl[3] br[3] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_6 
+ bl[4] br[4] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_7 
+ bl[5] br[5] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_8 
+ bl[6] br[6] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_9 
+ bl[7] br[7] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_10 
+ bl[8] br[8] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_11 
+ bl[9] br[9] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_12 
+ bl[10] br[10] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_13 
+ bl[11] br[11] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_14 
+ bl[12] br[12] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_15 
+ bl[13] br[13] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_16 
+ bl[14] br[14] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_17 
+ bl[15] br[15] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_18 
+ bl[16] br[16] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_19 
+ bl[17] br[17] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_20 
+ bl[18] br[18] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_21 
+ bl[19] br[19] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_22 
+ bl[20] br[20] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_23 
+ bl[21] br[21] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_24 
+ bl[22] br[22] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_25 
+ bl[23] br[23] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_26 
+ bl[24] br[24] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_27 
+ bl[25] br[25] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_28 
+ bl[26] br[26] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_29 
+ bl[27] br[27] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_30 
+ bl[28] br[28] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_31 
+ bl[29] br[29] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_32 
+ bl[30] br[30] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_33 
+ bl[31] br[31] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_34 
+ bl[32] br[32] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_35 
+ bl[33] br[33] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_36 
+ bl[34] br[34] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_37 
+ bl[35] br[35] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_38 
+ bl[36] br[36] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_39 
+ bl[37] br[37] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_40 
+ bl[38] br[38] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_41 
+ bl[39] br[39] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_42 
+ bl[40] br[40] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_43 
+ bl[41] br[41] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_44 
+ bl[42] br[42] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_45 
+ bl[43] br[43] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_46 
+ bl[44] br[44] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_47 
+ bl[45] br[45] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_48 
+ bl[46] br[46] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_49 
+ bl[47] br[47] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_50 
+ bl[48] br[48] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_51 
+ bl[49] br[49] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_52 
+ bl[50] br[50] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_53 
+ bl[51] br[51] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_54 
+ bl[52] br[52] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_55 
+ bl[53] br[53] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_56 
+ bl[54] br[54] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_57 
+ bl[55] br[55] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_58 
+ bl[56] br[56] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_59 
+ bl[57] br[57] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_60 
+ bl[58] br[58] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_61 
+ bl[59] br[59] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_62 
+ bl[60] br[60] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_63 
+ bl[61] br[61] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_64 
+ bl[62] br[62] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_65 
+ bl[63] br[63] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_66 
+ bl[64] br[64] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_67 
+ bl[65] br[65] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_68 
+ bl[66] br[66] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_69 
+ bl[67] br[67] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_70 
+ bl[68] br[68] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_71 
+ bl[69] br[69] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_72 
+ bl[70] br[70] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_73 
+ bl[71] br[71] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_74 
+ bl[72] br[72] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_75 
+ bl[73] br[73] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_76 
+ bl[74] br[74] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_77 
+ bl[75] br[75] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_78 
+ bl[76] br[76] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_79 
+ bl[77] br[77] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_80 
+ bl[78] br[78] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_81 
+ bl[79] br[79] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_82 
+ bl[80] br[80] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_83 
+ bl[81] br[81] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_84 
+ bl[82] br[82] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_85 
+ bl[83] br[83] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_86 
+ bl[84] br[84] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_87 
+ bl[85] br[85] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_88 
+ bl[86] br[86] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_89 
+ bl[87] br[87] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_90 
+ bl[88] br[88] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_91 
+ bl[89] br[89] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_92 
+ bl[90] br[90] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_93 
+ bl[91] br[91] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_94 
+ bl[92] br[92] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_95 
+ bl[93] br[93] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_96 
+ bl[94] br[94] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_97 
+ bl[95] br[95] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_98 
+ bl[96] br[96] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_99 
+ bl[97] br[97] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_100 
+ bl[98] br[98] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_101 
+ bl[99] br[99] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_102 
+ bl[100] br[100] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_103 
+ bl[101] br[101] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_104 
+ bl[102] br[102] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_105 
+ bl[103] br[103] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_106 
+ bl[104] br[104] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_107 
+ bl[105] br[105] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_108 
+ bl[106] br[106] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_109 
+ bl[107] br[107] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_110 
+ bl[108] br[108] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_111 
+ bl[109] br[109] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_112 
+ bl[110] br[110] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_113 
+ bl[111] br[111] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_114 
+ bl[112] br[112] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_115 
+ bl[113] br[113] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_116 
+ bl[114] br[114] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_117 
+ bl[115] br[115] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_118 
+ bl[116] br[116] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_119 
+ bl[117] br[117] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_120 
+ bl[118] br[118] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_121 
+ bl[119] br[119] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_122 
+ bl[120] br[120] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_123 
+ bl[121] br[121] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_124 
+ bl[122] br[122] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_125 
+ bl[123] br[123] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_126 
+ bl[124] br[124] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_127 
+ bl[125] br[125] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_128 
+ bl[126] br[126] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_129 
+ bl[127] br[127] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_130 
+ vdd vdd vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_131 
+ vdd vdd vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_0 
+ vdd vdd vss vdd vpb vnb wl[23] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_25_1 
+ rbl rbr vss vdd vpb vnb wl[23] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_25_2 
+ bl[0] br[0] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_3 
+ bl[1] br[1] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_4 
+ bl[2] br[2] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_5 
+ bl[3] br[3] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_6 
+ bl[4] br[4] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_7 
+ bl[5] br[5] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_8 
+ bl[6] br[6] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_9 
+ bl[7] br[7] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_10 
+ bl[8] br[8] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_11 
+ bl[9] br[9] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_12 
+ bl[10] br[10] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_13 
+ bl[11] br[11] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_14 
+ bl[12] br[12] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_15 
+ bl[13] br[13] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_16 
+ bl[14] br[14] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_17 
+ bl[15] br[15] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_18 
+ bl[16] br[16] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_19 
+ bl[17] br[17] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_20 
+ bl[18] br[18] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_21 
+ bl[19] br[19] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_22 
+ bl[20] br[20] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_23 
+ bl[21] br[21] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_24 
+ bl[22] br[22] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_25 
+ bl[23] br[23] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_26 
+ bl[24] br[24] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_27 
+ bl[25] br[25] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_28 
+ bl[26] br[26] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_29 
+ bl[27] br[27] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_30 
+ bl[28] br[28] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_31 
+ bl[29] br[29] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_32 
+ bl[30] br[30] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_33 
+ bl[31] br[31] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_34 
+ bl[32] br[32] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_35 
+ bl[33] br[33] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_36 
+ bl[34] br[34] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_37 
+ bl[35] br[35] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_38 
+ bl[36] br[36] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_39 
+ bl[37] br[37] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_40 
+ bl[38] br[38] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_41 
+ bl[39] br[39] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_42 
+ bl[40] br[40] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_43 
+ bl[41] br[41] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_44 
+ bl[42] br[42] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_45 
+ bl[43] br[43] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_46 
+ bl[44] br[44] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_47 
+ bl[45] br[45] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_48 
+ bl[46] br[46] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_49 
+ bl[47] br[47] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_50 
+ bl[48] br[48] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_51 
+ bl[49] br[49] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_52 
+ bl[50] br[50] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_53 
+ bl[51] br[51] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_54 
+ bl[52] br[52] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_55 
+ bl[53] br[53] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_56 
+ bl[54] br[54] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_57 
+ bl[55] br[55] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_58 
+ bl[56] br[56] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_59 
+ bl[57] br[57] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_60 
+ bl[58] br[58] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_61 
+ bl[59] br[59] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_62 
+ bl[60] br[60] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_63 
+ bl[61] br[61] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_64 
+ bl[62] br[62] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_65 
+ bl[63] br[63] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_66 
+ bl[64] br[64] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_67 
+ bl[65] br[65] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_68 
+ bl[66] br[66] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_69 
+ bl[67] br[67] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_70 
+ bl[68] br[68] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_71 
+ bl[69] br[69] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_72 
+ bl[70] br[70] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_73 
+ bl[71] br[71] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_74 
+ bl[72] br[72] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_75 
+ bl[73] br[73] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_76 
+ bl[74] br[74] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_77 
+ bl[75] br[75] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_78 
+ bl[76] br[76] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_79 
+ bl[77] br[77] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_80 
+ bl[78] br[78] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_81 
+ bl[79] br[79] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_82 
+ bl[80] br[80] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_83 
+ bl[81] br[81] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_84 
+ bl[82] br[82] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_85 
+ bl[83] br[83] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_86 
+ bl[84] br[84] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_87 
+ bl[85] br[85] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_88 
+ bl[86] br[86] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_89 
+ bl[87] br[87] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_90 
+ bl[88] br[88] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_91 
+ bl[89] br[89] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_92 
+ bl[90] br[90] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_93 
+ bl[91] br[91] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_94 
+ bl[92] br[92] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_95 
+ bl[93] br[93] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_96 
+ bl[94] br[94] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_97 
+ bl[95] br[95] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_98 
+ bl[96] br[96] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_99 
+ bl[97] br[97] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_100 
+ bl[98] br[98] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_101 
+ bl[99] br[99] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_102 
+ bl[100] br[100] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_103 
+ bl[101] br[101] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_104 
+ bl[102] br[102] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_105 
+ bl[103] br[103] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_106 
+ bl[104] br[104] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_107 
+ bl[105] br[105] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_108 
+ bl[106] br[106] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_109 
+ bl[107] br[107] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_110 
+ bl[108] br[108] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_111 
+ bl[109] br[109] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_112 
+ bl[110] br[110] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_113 
+ bl[111] br[111] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_114 
+ bl[112] br[112] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_115 
+ bl[113] br[113] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_116 
+ bl[114] br[114] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_117 
+ bl[115] br[115] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_118 
+ bl[116] br[116] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_119 
+ bl[117] br[117] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_120 
+ bl[118] br[118] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_121 
+ bl[119] br[119] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_122 
+ bl[120] br[120] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_123 
+ bl[121] br[121] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_124 
+ bl[122] br[122] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_125 
+ bl[123] br[123] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_126 
+ bl[124] br[124] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_127 
+ bl[125] br[125] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_128 
+ bl[126] br[126] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_129 
+ bl[127] br[127] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_130 
+ vdd vdd vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_131 
+ vdd vdd vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_0 
+ vdd vdd vss vdd vpb vnb wl[24] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_26_1 
+ rbl rbr vss vdd vpb vnb wl[24] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_26_2 
+ bl[0] br[0] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_3 
+ bl[1] br[1] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_4 
+ bl[2] br[2] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_5 
+ bl[3] br[3] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_6 
+ bl[4] br[4] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_7 
+ bl[5] br[5] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_8 
+ bl[6] br[6] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_9 
+ bl[7] br[7] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_10 
+ bl[8] br[8] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_11 
+ bl[9] br[9] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_12 
+ bl[10] br[10] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_13 
+ bl[11] br[11] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_14 
+ bl[12] br[12] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_15 
+ bl[13] br[13] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_16 
+ bl[14] br[14] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_17 
+ bl[15] br[15] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_18 
+ bl[16] br[16] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_19 
+ bl[17] br[17] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_20 
+ bl[18] br[18] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_21 
+ bl[19] br[19] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_22 
+ bl[20] br[20] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_23 
+ bl[21] br[21] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_24 
+ bl[22] br[22] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_25 
+ bl[23] br[23] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_26 
+ bl[24] br[24] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_27 
+ bl[25] br[25] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_28 
+ bl[26] br[26] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_29 
+ bl[27] br[27] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_30 
+ bl[28] br[28] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_31 
+ bl[29] br[29] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_32 
+ bl[30] br[30] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_33 
+ bl[31] br[31] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_34 
+ bl[32] br[32] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_35 
+ bl[33] br[33] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_36 
+ bl[34] br[34] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_37 
+ bl[35] br[35] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_38 
+ bl[36] br[36] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_39 
+ bl[37] br[37] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_40 
+ bl[38] br[38] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_41 
+ bl[39] br[39] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_42 
+ bl[40] br[40] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_43 
+ bl[41] br[41] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_44 
+ bl[42] br[42] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_45 
+ bl[43] br[43] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_46 
+ bl[44] br[44] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_47 
+ bl[45] br[45] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_48 
+ bl[46] br[46] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_49 
+ bl[47] br[47] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_50 
+ bl[48] br[48] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_51 
+ bl[49] br[49] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_52 
+ bl[50] br[50] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_53 
+ bl[51] br[51] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_54 
+ bl[52] br[52] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_55 
+ bl[53] br[53] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_56 
+ bl[54] br[54] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_57 
+ bl[55] br[55] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_58 
+ bl[56] br[56] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_59 
+ bl[57] br[57] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_60 
+ bl[58] br[58] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_61 
+ bl[59] br[59] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_62 
+ bl[60] br[60] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_63 
+ bl[61] br[61] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_64 
+ bl[62] br[62] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_65 
+ bl[63] br[63] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_66 
+ bl[64] br[64] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_67 
+ bl[65] br[65] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_68 
+ bl[66] br[66] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_69 
+ bl[67] br[67] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_70 
+ bl[68] br[68] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_71 
+ bl[69] br[69] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_72 
+ bl[70] br[70] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_73 
+ bl[71] br[71] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_74 
+ bl[72] br[72] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_75 
+ bl[73] br[73] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_76 
+ bl[74] br[74] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_77 
+ bl[75] br[75] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_78 
+ bl[76] br[76] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_79 
+ bl[77] br[77] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_80 
+ bl[78] br[78] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_81 
+ bl[79] br[79] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_82 
+ bl[80] br[80] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_83 
+ bl[81] br[81] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_84 
+ bl[82] br[82] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_85 
+ bl[83] br[83] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_86 
+ bl[84] br[84] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_87 
+ bl[85] br[85] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_88 
+ bl[86] br[86] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_89 
+ bl[87] br[87] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_90 
+ bl[88] br[88] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_91 
+ bl[89] br[89] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_92 
+ bl[90] br[90] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_93 
+ bl[91] br[91] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_94 
+ bl[92] br[92] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_95 
+ bl[93] br[93] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_96 
+ bl[94] br[94] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_97 
+ bl[95] br[95] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_98 
+ bl[96] br[96] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_99 
+ bl[97] br[97] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_100 
+ bl[98] br[98] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_101 
+ bl[99] br[99] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_102 
+ bl[100] br[100] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_103 
+ bl[101] br[101] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_104 
+ bl[102] br[102] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_105 
+ bl[103] br[103] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_106 
+ bl[104] br[104] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_107 
+ bl[105] br[105] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_108 
+ bl[106] br[106] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_109 
+ bl[107] br[107] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_110 
+ bl[108] br[108] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_111 
+ bl[109] br[109] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_112 
+ bl[110] br[110] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_113 
+ bl[111] br[111] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_114 
+ bl[112] br[112] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_115 
+ bl[113] br[113] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_116 
+ bl[114] br[114] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_117 
+ bl[115] br[115] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_118 
+ bl[116] br[116] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_119 
+ bl[117] br[117] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_120 
+ bl[118] br[118] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_121 
+ bl[119] br[119] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_122 
+ bl[120] br[120] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_123 
+ bl[121] br[121] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_124 
+ bl[122] br[122] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_125 
+ bl[123] br[123] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_126 
+ bl[124] br[124] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_127 
+ bl[125] br[125] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_128 
+ bl[126] br[126] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_129 
+ bl[127] br[127] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_130 
+ vdd vdd vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_131 
+ vdd vdd vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_0 
+ vdd vdd vss vdd vpb vnb wl[25] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_27_1 
+ rbl rbr vss vdd vpb vnb wl[25] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_27_2 
+ bl[0] br[0] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_3 
+ bl[1] br[1] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_4 
+ bl[2] br[2] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_5 
+ bl[3] br[3] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_6 
+ bl[4] br[4] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_7 
+ bl[5] br[5] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_8 
+ bl[6] br[6] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_9 
+ bl[7] br[7] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_10 
+ bl[8] br[8] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_11 
+ bl[9] br[9] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_12 
+ bl[10] br[10] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_13 
+ bl[11] br[11] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_14 
+ bl[12] br[12] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_15 
+ bl[13] br[13] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_16 
+ bl[14] br[14] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_17 
+ bl[15] br[15] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_18 
+ bl[16] br[16] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_19 
+ bl[17] br[17] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_20 
+ bl[18] br[18] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_21 
+ bl[19] br[19] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_22 
+ bl[20] br[20] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_23 
+ bl[21] br[21] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_24 
+ bl[22] br[22] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_25 
+ bl[23] br[23] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_26 
+ bl[24] br[24] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_27 
+ bl[25] br[25] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_28 
+ bl[26] br[26] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_29 
+ bl[27] br[27] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_30 
+ bl[28] br[28] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_31 
+ bl[29] br[29] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_32 
+ bl[30] br[30] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_33 
+ bl[31] br[31] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_34 
+ bl[32] br[32] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_35 
+ bl[33] br[33] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_36 
+ bl[34] br[34] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_37 
+ bl[35] br[35] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_38 
+ bl[36] br[36] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_39 
+ bl[37] br[37] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_40 
+ bl[38] br[38] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_41 
+ bl[39] br[39] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_42 
+ bl[40] br[40] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_43 
+ bl[41] br[41] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_44 
+ bl[42] br[42] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_45 
+ bl[43] br[43] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_46 
+ bl[44] br[44] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_47 
+ bl[45] br[45] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_48 
+ bl[46] br[46] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_49 
+ bl[47] br[47] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_50 
+ bl[48] br[48] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_51 
+ bl[49] br[49] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_52 
+ bl[50] br[50] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_53 
+ bl[51] br[51] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_54 
+ bl[52] br[52] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_55 
+ bl[53] br[53] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_56 
+ bl[54] br[54] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_57 
+ bl[55] br[55] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_58 
+ bl[56] br[56] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_59 
+ bl[57] br[57] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_60 
+ bl[58] br[58] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_61 
+ bl[59] br[59] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_62 
+ bl[60] br[60] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_63 
+ bl[61] br[61] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_64 
+ bl[62] br[62] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_65 
+ bl[63] br[63] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_66 
+ bl[64] br[64] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_67 
+ bl[65] br[65] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_68 
+ bl[66] br[66] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_69 
+ bl[67] br[67] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_70 
+ bl[68] br[68] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_71 
+ bl[69] br[69] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_72 
+ bl[70] br[70] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_73 
+ bl[71] br[71] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_74 
+ bl[72] br[72] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_75 
+ bl[73] br[73] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_76 
+ bl[74] br[74] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_77 
+ bl[75] br[75] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_78 
+ bl[76] br[76] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_79 
+ bl[77] br[77] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_80 
+ bl[78] br[78] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_81 
+ bl[79] br[79] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_82 
+ bl[80] br[80] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_83 
+ bl[81] br[81] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_84 
+ bl[82] br[82] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_85 
+ bl[83] br[83] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_86 
+ bl[84] br[84] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_87 
+ bl[85] br[85] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_88 
+ bl[86] br[86] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_89 
+ bl[87] br[87] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_90 
+ bl[88] br[88] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_91 
+ bl[89] br[89] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_92 
+ bl[90] br[90] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_93 
+ bl[91] br[91] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_94 
+ bl[92] br[92] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_95 
+ bl[93] br[93] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_96 
+ bl[94] br[94] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_97 
+ bl[95] br[95] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_98 
+ bl[96] br[96] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_99 
+ bl[97] br[97] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_100 
+ bl[98] br[98] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_101 
+ bl[99] br[99] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_102 
+ bl[100] br[100] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_103 
+ bl[101] br[101] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_104 
+ bl[102] br[102] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_105 
+ bl[103] br[103] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_106 
+ bl[104] br[104] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_107 
+ bl[105] br[105] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_108 
+ bl[106] br[106] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_109 
+ bl[107] br[107] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_110 
+ bl[108] br[108] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_111 
+ bl[109] br[109] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_112 
+ bl[110] br[110] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_113 
+ bl[111] br[111] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_114 
+ bl[112] br[112] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_115 
+ bl[113] br[113] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_116 
+ bl[114] br[114] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_117 
+ bl[115] br[115] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_118 
+ bl[116] br[116] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_119 
+ bl[117] br[117] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_120 
+ bl[118] br[118] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_121 
+ bl[119] br[119] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_122 
+ bl[120] br[120] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_123 
+ bl[121] br[121] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_124 
+ bl[122] br[122] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_125 
+ bl[123] br[123] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_126 
+ bl[124] br[124] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_127 
+ bl[125] br[125] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_128 
+ bl[126] br[126] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_129 
+ bl[127] br[127] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_130 
+ vdd vdd vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_131 
+ vdd vdd vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_0 
+ vdd vdd vss vdd vpb vnb wl[26] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_28_1 
+ rbl rbr vss vdd vpb vnb wl[26] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_28_2 
+ bl[0] br[0] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_3 
+ bl[1] br[1] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_4 
+ bl[2] br[2] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_5 
+ bl[3] br[3] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_6 
+ bl[4] br[4] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_7 
+ bl[5] br[5] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_8 
+ bl[6] br[6] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_9 
+ bl[7] br[7] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_10 
+ bl[8] br[8] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_11 
+ bl[9] br[9] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_12 
+ bl[10] br[10] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_13 
+ bl[11] br[11] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_14 
+ bl[12] br[12] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_15 
+ bl[13] br[13] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_16 
+ bl[14] br[14] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_17 
+ bl[15] br[15] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_18 
+ bl[16] br[16] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_19 
+ bl[17] br[17] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_20 
+ bl[18] br[18] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_21 
+ bl[19] br[19] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_22 
+ bl[20] br[20] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_23 
+ bl[21] br[21] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_24 
+ bl[22] br[22] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_25 
+ bl[23] br[23] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_26 
+ bl[24] br[24] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_27 
+ bl[25] br[25] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_28 
+ bl[26] br[26] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_29 
+ bl[27] br[27] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_30 
+ bl[28] br[28] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_31 
+ bl[29] br[29] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_32 
+ bl[30] br[30] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_33 
+ bl[31] br[31] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_34 
+ bl[32] br[32] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_35 
+ bl[33] br[33] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_36 
+ bl[34] br[34] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_37 
+ bl[35] br[35] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_38 
+ bl[36] br[36] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_39 
+ bl[37] br[37] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_40 
+ bl[38] br[38] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_41 
+ bl[39] br[39] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_42 
+ bl[40] br[40] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_43 
+ bl[41] br[41] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_44 
+ bl[42] br[42] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_45 
+ bl[43] br[43] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_46 
+ bl[44] br[44] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_47 
+ bl[45] br[45] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_48 
+ bl[46] br[46] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_49 
+ bl[47] br[47] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_50 
+ bl[48] br[48] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_51 
+ bl[49] br[49] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_52 
+ bl[50] br[50] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_53 
+ bl[51] br[51] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_54 
+ bl[52] br[52] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_55 
+ bl[53] br[53] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_56 
+ bl[54] br[54] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_57 
+ bl[55] br[55] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_58 
+ bl[56] br[56] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_59 
+ bl[57] br[57] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_60 
+ bl[58] br[58] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_61 
+ bl[59] br[59] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_62 
+ bl[60] br[60] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_63 
+ bl[61] br[61] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_64 
+ bl[62] br[62] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_65 
+ bl[63] br[63] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_66 
+ bl[64] br[64] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_67 
+ bl[65] br[65] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_68 
+ bl[66] br[66] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_69 
+ bl[67] br[67] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_70 
+ bl[68] br[68] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_71 
+ bl[69] br[69] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_72 
+ bl[70] br[70] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_73 
+ bl[71] br[71] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_74 
+ bl[72] br[72] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_75 
+ bl[73] br[73] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_76 
+ bl[74] br[74] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_77 
+ bl[75] br[75] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_78 
+ bl[76] br[76] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_79 
+ bl[77] br[77] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_80 
+ bl[78] br[78] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_81 
+ bl[79] br[79] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_82 
+ bl[80] br[80] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_83 
+ bl[81] br[81] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_84 
+ bl[82] br[82] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_85 
+ bl[83] br[83] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_86 
+ bl[84] br[84] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_87 
+ bl[85] br[85] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_88 
+ bl[86] br[86] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_89 
+ bl[87] br[87] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_90 
+ bl[88] br[88] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_91 
+ bl[89] br[89] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_92 
+ bl[90] br[90] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_93 
+ bl[91] br[91] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_94 
+ bl[92] br[92] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_95 
+ bl[93] br[93] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_96 
+ bl[94] br[94] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_97 
+ bl[95] br[95] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_98 
+ bl[96] br[96] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_99 
+ bl[97] br[97] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_100 
+ bl[98] br[98] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_101 
+ bl[99] br[99] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_102 
+ bl[100] br[100] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_103 
+ bl[101] br[101] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_104 
+ bl[102] br[102] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_105 
+ bl[103] br[103] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_106 
+ bl[104] br[104] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_107 
+ bl[105] br[105] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_108 
+ bl[106] br[106] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_109 
+ bl[107] br[107] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_110 
+ bl[108] br[108] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_111 
+ bl[109] br[109] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_112 
+ bl[110] br[110] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_113 
+ bl[111] br[111] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_114 
+ bl[112] br[112] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_115 
+ bl[113] br[113] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_116 
+ bl[114] br[114] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_117 
+ bl[115] br[115] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_118 
+ bl[116] br[116] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_119 
+ bl[117] br[117] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_120 
+ bl[118] br[118] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_121 
+ bl[119] br[119] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_122 
+ bl[120] br[120] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_123 
+ bl[121] br[121] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_124 
+ bl[122] br[122] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_125 
+ bl[123] br[123] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_126 
+ bl[124] br[124] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_127 
+ bl[125] br[125] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_128 
+ bl[126] br[126] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_129 
+ bl[127] br[127] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_130 
+ vdd vdd vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_131 
+ vdd vdd vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_0 
+ vdd vdd vss vdd vpb vnb wl[27] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_29_1 
+ rbl rbr vss vdd vpb vnb wl[27] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_29_2 
+ bl[0] br[0] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_3 
+ bl[1] br[1] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_4 
+ bl[2] br[2] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_5 
+ bl[3] br[3] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_6 
+ bl[4] br[4] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_7 
+ bl[5] br[5] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_8 
+ bl[6] br[6] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_9 
+ bl[7] br[7] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_10 
+ bl[8] br[8] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_11 
+ bl[9] br[9] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_12 
+ bl[10] br[10] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_13 
+ bl[11] br[11] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_14 
+ bl[12] br[12] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_15 
+ bl[13] br[13] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_16 
+ bl[14] br[14] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_17 
+ bl[15] br[15] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_18 
+ bl[16] br[16] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_19 
+ bl[17] br[17] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_20 
+ bl[18] br[18] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_21 
+ bl[19] br[19] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_22 
+ bl[20] br[20] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_23 
+ bl[21] br[21] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_24 
+ bl[22] br[22] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_25 
+ bl[23] br[23] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_26 
+ bl[24] br[24] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_27 
+ bl[25] br[25] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_28 
+ bl[26] br[26] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_29 
+ bl[27] br[27] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_30 
+ bl[28] br[28] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_31 
+ bl[29] br[29] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_32 
+ bl[30] br[30] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_33 
+ bl[31] br[31] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_34 
+ bl[32] br[32] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_35 
+ bl[33] br[33] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_36 
+ bl[34] br[34] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_37 
+ bl[35] br[35] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_38 
+ bl[36] br[36] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_39 
+ bl[37] br[37] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_40 
+ bl[38] br[38] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_41 
+ bl[39] br[39] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_42 
+ bl[40] br[40] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_43 
+ bl[41] br[41] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_44 
+ bl[42] br[42] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_45 
+ bl[43] br[43] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_46 
+ bl[44] br[44] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_47 
+ bl[45] br[45] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_48 
+ bl[46] br[46] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_49 
+ bl[47] br[47] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_50 
+ bl[48] br[48] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_51 
+ bl[49] br[49] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_52 
+ bl[50] br[50] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_53 
+ bl[51] br[51] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_54 
+ bl[52] br[52] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_55 
+ bl[53] br[53] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_56 
+ bl[54] br[54] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_57 
+ bl[55] br[55] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_58 
+ bl[56] br[56] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_59 
+ bl[57] br[57] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_60 
+ bl[58] br[58] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_61 
+ bl[59] br[59] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_62 
+ bl[60] br[60] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_63 
+ bl[61] br[61] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_64 
+ bl[62] br[62] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_65 
+ bl[63] br[63] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_66 
+ bl[64] br[64] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_67 
+ bl[65] br[65] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_68 
+ bl[66] br[66] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_69 
+ bl[67] br[67] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_70 
+ bl[68] br[68] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_71 
+ bl[69] br[69] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_72 
+ bl[70] br[70] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_73 
+ bl[71] br[71] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_74 
+ bl[72] br[72] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_75 
+ bl[73] br[73] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_76 
+ bl[74] br[74] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_77 
+ bl[75] br[75] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_78 
+ bl[76] br[76] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_79 
+ bl[77] br[77] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_80 
+ bl[78] br[78] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_81 
+ bl[79] br[79] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_82 
+ bl[80] br[80] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_83 
+ bl[81] br[81] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_84 
+ bl[82] br[82] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_85 
+ bl[83] br[83] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_86 
+ bl[84] br[84] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_87 
+ bl[85] br[85] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_88 
+ bl[86] br[86] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_89 
+ bl[87] br[87] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_90 
+ bl[88] br[88] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_91 
+ bl[89] br[89] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_92 
+ bl[90] br[90] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_93 
+ bl[91] br[91] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_94 
+ bl[92] br[92] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_95 
+ bl[93] br[93] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_96 
+ bl[94] br[94] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_97 
+ bl[95] br[95] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_98 
+ bl[96] br[96] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_99 
+ bl[97] br[97] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_100 
+ bl[98] br[98] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_101 
+ bl[99] br[99] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_102 
+ bl[100] br[100] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_103 
+ bl[101] br[101] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_104 
+ bl[102] br[102] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_105 
+ bl[103] br[103] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_106 
+ bl[104] br[104] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_107 
+ bl[105] br[105] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_108 
+ bl[106] br[106] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_109 
+ bl[107] br[107] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_110 
+ bl[108] br[108] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_111 
+ bl[109] br[109] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_112 
+ bl[110] br[110] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_113 
+ bl[111] br[111] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_114 
+ bl[112] br[112] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_115 
+ bl[113] br[113] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_116 
+ bl[114] br[114] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_117 
+ bl[115] br[115] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_118 
+ bl[116] br[116] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_119 
+ bl[117] br[117] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_120 
+ bl[118] br[118] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_121 
+ bl[119] br[119] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_122 
+ bl[120] br[120] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_123 
+ bl[121] br[121] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_124 
+ bl[122] br[122] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_125 
+ bl[123] br[123] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_126 
+ bl[124] br[124] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_127 
+ bl[125] br[125] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_128 
+ bl[126] br[126] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_129 
+ bl[127] br[127] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_130 
+ vdd vdd vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_131 
+ vdd vdd vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_0 
+ vdd vdd vss vdd vpb vnb wl[28] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_30_1 
+ rbl rbr vss vdd vpb vnb wl[28] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_30_2 
+ bl[0] br[0] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_3 
+ bl[1] br[1] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_4 
+ bl[2] br[2] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_5 
+ bl[3] br[3] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_6 
+ bl[4] br[4] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_7 
+ bl[5] br[5] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_8 
+ bl[6] br[6] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_9 
+ bl[7] br[7] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_10 
+ bl[8] br[8] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_11 
+ bl[9] br[9] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_12 
+ bl[10] br[10] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_13 
+ bl[11] br[11] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_14 
+ bl[12] br[12] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_15 
+ bl[13] br[13] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_16 
+ bl[14] br[14] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_17 
+ bl[15] br[15] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_18 
+ bl[16] br[16] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_19 
+ bl[17] br[17] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_20 
+ bl[18] br[18] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_21 
+ bl[19] br[19] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_22 
+ bl[20] br[20] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_23 
+ bl[21] br[21] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_24 
+ bl[22] br[22] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_25 
+ bl[23] br[23] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_26 
+ bl[24] br[24] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_27 
+ bl[25] br[25] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_28 
+ bl[26] br[26] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_29 
+ bl[27] br[27] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_30 
+ bl[28] br[28] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_31 
+ bl[29] br[29] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_32 
+ bl[30] br[30] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_33 
+ bl[31] br[31] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_34 
+ bl[32] br[32] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_35 
+ bl[33] br[33] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_36 
+ bl[34] br[34] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_37 
+ bl[35] br[35] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_38 
+ bl[36] br[36] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_39 
+ bl[37] br[37] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_40 
+ bl[38] br[38] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_41 
+ bl[39] br[39] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_42 
+ bl[40] br[40] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_43 
+ bl[41] br[41] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_44 
+ bl[42] br[42] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_45 
+ bl[43] br[43] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_46 
+ bl[44] br[44] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_47 
+ bl[45] br[45] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_48 
+ bl[46] br[46] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_49 
+ bl[47] br[47] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_50 
+ bl[48] br[48] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_51 
+ bl[49] br[49] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_52 
+ bl[50] br[50] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_53 
+ bl[51] br[51] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_54 
+ bl[52] br[52] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_55 
+ bl[53] br[53] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_56 
+ bl[54] br[54] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_57 
+ bl[55] br[55] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_58 
+ bl[56] br[56] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_59 
+ bl[57] br[57] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_60 
+ bl[58] br[58] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_61 
+ bl[59] br[59] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_62 
+ bl[60] br[60] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_63 
+ bl[61] br[61] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_64 
+ bl[62] br[62] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_65 
+ bl[63] br[63] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_66 
+ bl[64] br[64] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_67 
+ bl[65] br[65] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_68 
+ bl[66] br[66] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_69 
+ bl[67] br[67] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_70 
+ bl[68] br[68] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_71 
+ bl[69] br[69] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_72 
+ bl[70] br[70] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_73 
+ bl[71] br[71] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_74 
+ bl[72] br[72] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_75 
+ bl[73] br[73] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_76 
+ bl[74] br[74] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_77 
+ bl[75] br[75] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_78 
+ bl[76] br[76] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_79 
+ bl[77] br[77] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_80 
+ bl[78] br[78] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_81 
+ bl[79] br[79] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_82 
+ bl[80] br[80] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_83 
+ bl[81] br[81] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_84 
+ bl[82] br[82] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_85 
+ bl[83] br[83] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_86 
+ bl[84] br[84] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_87 
+ bl[85] br[85] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_88 
+ bl[86] br[86] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_89 
+ bl[87] br[87] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_90 
+ bl[88] br[88] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_91 
+ bl[89] br[89] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_92 
+ bl[90] br[90] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_93 
+ bl[91] br[91] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_94 
+ bl[92] br[92] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_95 
+ bl[93] br[93] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_96 
+ bl[94] br[94] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_97 
+ bl[95] br[95] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_98 
+ bl[96] br[96] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_99 
+ bl[97] br[97] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_100 
+ bl[98] br[98] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_101 
+ bl[99] br[99] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_102 
+ bl[100] br[100] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_103 
+ bl[101] br[101] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_104 
+ bl[102] br[102] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_105 
+ bl[103] br[103] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_106 
+ bl[104] br[104] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_107 
+ bl[105] br[105] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_108 
+ bl[106] br[106] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_109 
+ bl[107] br[107] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_110 
+ bl[108] br[108] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_111 
+ bl[109] br[109] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_112 
+ bl[110] br[110] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_113 
+ bl[111] br[111] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_114 
+ bl[112] br[112] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_115 
+ bl[113] br[113] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_116 
+ bl[114] br[114] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_117 
+ bl[115] br[115] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_118 
+ bl[116] br[116] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_119 
+ bl[117] br[117] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_120 
+ bl[118] br[118] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_121 
+ bl[119] br[119] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_122 
+ bl[120] br[120] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_123 
+ bl[121] br[121] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_124 
+ bl[122] br[122] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_125 
+ bl[123] br[123] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_126 
+ bl[124] br[124] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_127 
+ bl[125] br[125] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_128 
+ bl[126] br[126] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_129 
+ bl[127] br[127] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_130 
+ vdd vdd vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_131 
+ vdd vdd vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_0 
+ vdd vdd vss vdd vpb vnb wl[29] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_31_1 
+ rbl rbr vss vdd vpb vnb wl[29] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_31_2 
+ bl[0] br[0] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_3 
+ bl[1] br[1] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_4 
+ bl[2] br[2] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_5 
+ bl[3] br[3] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_6 
+ bl[4] br[4] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_7 
+ bl[5] br[5] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_8 
+ bl[6] br[6] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_9 
+ bl[7] br[7] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_10 
+ bl[8] br[8] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_11 
+ bl[9] br[9] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_12 
+ bl[10] br[10] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_13 
+ bl[11] br[11] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_14 
+ bl[12] br[12] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_15 
+ bl[13] br[13] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_16 
+ bl[14] br[14] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_17 
+ bl[15] br[15] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_18 
+ bl[16] br[16] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_19 
+ bl[17] br[17] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_20 
+ bl[18] br[18] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_21 
+ bl[19] br[19] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_22 
+ bl[20] br[20] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_23 
+ bl[21] br[21] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_24 
+ bl[22] br[22] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_25 
+ bl[23] br[23] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_26 
+ bl[24] br[24] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_27 
+ bl[25] br[25] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_28 
+ bl[26] br[26] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_29 
+ bl[27] br[27] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_30 
+ bl[28] br[28] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_31 
+ bl[29] br[29] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_32 
+ bl[30] br[30] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_33 
+ bl[31] br[31] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_34 
+ bl[32] br[32] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_35 
+ bl[33] br[33] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_36 
+ bl[34] br[34] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_37 
+ bl[35] br[35] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_38 
+ bl[36] br[36] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_39 
+ bl[37] br[37] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_40 
+ bl[38] br[38] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_41 
+ bl[39] br[39] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_42 
+ bl[40] br[40] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_43 
+ bl[41] br[41] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_44 
+ bl[42] br[42] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_45 
+ bl[43] br[43] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_46 
+ bl[44] br[44] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_47 
+ bl[45] br[45] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_48 
+ bl[46] br[46] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_49 
+ bl[47] br[47] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_50 
+ bl[48] br[48] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_51 
+ bl[49] br[49] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_52 
+ bl[50] br[50] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_53 
+ bl[51] br[51] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_54 
+ bl[52] br[52] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_55 
+ bl[53] br[53] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_56 
+ bl[54] br[54] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_57 
+ bl[55] br[55] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_58 
+ bl[56] br[56] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_59 
+ bl[57] br[57] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_60 
+ bl[58] br[58] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_61 
+ bl[59] br[59] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_62 
+ bl[60] br[60] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_63 
+ bl[61] br[61] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_64 
+ bl[62] br[62] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_65 
+ bl[63] br[63] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_66 
+ bl[64] br[64] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_67 
+ bl[65] br[65] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_68 
+ bl[66] br[66] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_69 
+ bl[67] br[67] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_70 
+ bl[68] br[68] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_71 
+ bl[69] br[69] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_72 
+ bl[70] br[70] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_73 
+ bl[71] br[71] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_74 
+ bl[72] br[72] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_75 
+ bl[73] br[73] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_76 
+ bl[74] br[74] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_77 
+ bl[75] br[75] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_78 
+ bl[76] br[76] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_79 
+ bl[77] br[77] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_80 
+ bl[78] br[78] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_81 
+ bl[79] br[79] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_82 
+ bl[80] br[80] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_83 
+ bl[81] br[81] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_84 
+ bl[82] br[82] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_85 
+ bl[83] br[83] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_86 
+ bl[84] br[84] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_87 
+ bl[85] br[85] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_88 
+ bl[86] br[86] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_89 
+ bl[87] br[87] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_90 
+ bl[88] br[88] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_91 
+ bl[89] br[89] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_92 
+ bl[90] br[90] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_93 
+ bl[91] br[91] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_94 
+ bl[92] br[92] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_95 
+ bl[93] br[93] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_96 
+ bl[94] br[94] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_97 
+ bl[95] br[95] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_98 
+ bl[96] br[96] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_99 
+ bl[97] br[97] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_100 
+ bl[98] br[98] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_101 
+ bl[99] br[99] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_102 
+ bl[100] br[100] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_103 
+ bl[101] br[101] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_104 
+ bl[102] br[102] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_105 
+ bl[103] br[103] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_106 
+ bl[104] br[104] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_107 
+ bl[105] br[105] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_108 
+ bl[106] br[106] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_109 
+ bl[107] br[107] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_110 
+ bl[108] br[108] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_111 
+ bl[109] br[109] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_112 
+ bl[110] br[110] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_113 
+ bl[111] br[111] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_114 
+ bl[112] br[112] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_115 
+ bl[113] br[113] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_116 
+ bl[114] br[114] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_117 
+ bl[115] br[115] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_118 
+ bl[116] br[116] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_119 
+ bl[117] br[117] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_120 
+ bl[118] br[118] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_121 
+ bl[119] br[119] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_122 
+ bl[120] br[120] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_123 
+ bl[121] br[121] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_124 
+ bl[122] br[122] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_125 
+ bl[123] br[123] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_126 
+ bl[124] br[124] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_127 
+ bl[125] br[125] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_128 
+ bl[126] br[126] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_129 
+ bl[127] br[127] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_130 
+ vdd vdd vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_131 
+ vdd vdd vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_0 
+ vdd vdd vss vdd vpb vnb wl[30] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_32_1 
+ rbl rbr vss vdd vpb vnb wl[30] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_32_2 
+ bl[0] br[0] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_3 
+ bl[1] br[1] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_4 
+ bl[2] br[2] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_5 
+ bl[3] br[3] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_6 
+ bl[4] br[4] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_7 
+ bl[5] br[5] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_8 
+ bl[6] br[6] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_9 
+ bl[7] br[7] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_10 
+ bl[8] br[8] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_11 
+ bl[9] br[9] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_12 
+ bl[10] br[10] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_13 
+ bl[11] br[11] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_14 
+ bl[12] br[12] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_15 
+ bl[13] br[13] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_16 
+ bl[14] br[14] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_17 
+ bl[15] br[15] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_18 
+ bl[16] br[16] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_19 
+ bl[17] br[17] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_20 
+ bl[18] br[18] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_21 
+ bl[19] br[19] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_22 
+ bl[20] br[20] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_23 
+ bl[21] br[21] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_24 
+ bl[22] br[22] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_25 
+ bl[23] br[23] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_26 
+ bl[24] br[24] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_27 
+ bl[25] br[25] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_28 
+ bl[26] br[26] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_29 
+ bl[27] br[27] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_30 
+ bl[28] br[28] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_31 
+ bl[29] br[29] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_32 
+ bl[30] br[30] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_33 
+ bl[31] br[31] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_34 
+ bl[32] br[32] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_35 
+ bl[33] br[33] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_36 
+ bl[34] br[34] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_37 
+ bl[35] br[35] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_38 
+ bl[36] br[36] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_39 
+ bl[37] br[37] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_40 
+ bl[38] br[38] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_41 
+ bl[39] br[39] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_42 
+ bl[40] br[40] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_43 
+ bl[41] br[41] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_44 
+ bl[42] br[42] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_45 
+ bl[43] br[43] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_46 
+ bl[44] br[44] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_47 
+ bl[45] br[45] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_48 
+ bl[46] br[46] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_49 
+ bl[47] br[47] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_50 
+ bl[48] br[48] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_51 
+ bl[49] br[49] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_52 
+ bl[50] br[50] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_53 
+ bl[51] br[51] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_54 
+ bl[52] br[52] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_55 
+ bl[53] br[53] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_56 
+ bl[54] br[54] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_57 
+ bl[55] br[55] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_58 
+ bl[56] br[56] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_59 
+ bl[57] br[57] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_60 
+ bl[58] br[58] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_61 
+ bl[59] br[59] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_62 
+ bl[60] br[60] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_63 
+ bl[61] br[61] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_64 
+ bl[62] br[62] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_65 
+ bl[63] br[63] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_66 
+ bl[64] br[64] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_67 
+ bl[65] br[65] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_68 
+ bl[66] br[66] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_69 
+ bl[67] br[67] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_70 
+ bl[68] br[68] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_71 
+ bl[69] br[69] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_72 
+ bl[70] br[70] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_73 
+ bl[71] br[71] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_74 
+ bl[72] br[72] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_75 
+ bl[73] br[73] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_76 
+ bl[74] br[74] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_77 
+ bl[75] br[75] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_78 
+ bl[76] br[76] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_79 
+ bl[77] br[77] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_80 
+ bl[78] br[78] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_81 
+ bl[79] br[79] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_82 
+ bl[80] br[80] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_83 
+ bl[81] br[81] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_84 
+ bl[82] br[82] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_85 
+ bl[83] br[83] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_86 
+ bl[84] br[84] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_87 
+ bl[85] br[85] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_88 
+ bl[86] br[86] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_89 
+ bl[87] br[87] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_90 
+ bl[88] br[88] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_91 
+ bl[89] br[89] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_92 
+ bl[90] br[90] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_93 
+ bl[91] br[91] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_94 
+ bl[92] br[92] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_95 
+ bl[93] br[93] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_96 
+ bl[94] br[94] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_97 
+ bl[95] br[95] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_98 
+ bl[96] br[96] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_99 
+ bl[97] br[97] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_100 
+ bl[98] br[98] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_101 
+ bl[99] br[99] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_102 
+ bl[100] br[100] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_103 
+ bl[101] br[101] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_104 
+ bl[102] br[102] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_105 
+ bl[103] br[103] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_106 
+ bl[104] br[104] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_107 
+ bl[105] br[105] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_108 
+ bl[106] br[106] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_109 
+ bl[107] br[107] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_110 
+ bl[108] br[108] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_111 
+ bl[109] br[109] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_112 
+ bl[110] br[110] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_113 
+ bl[111] br[111] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_114 
+ bl[112] br[112] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_115 
+ bl[113] br[113] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_116 
+ bl[114] br[114] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_117 
+ bl[115] br[115] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_118 
+ bl[116] br[116] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_119 
+ bl[117] br[117] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_120 
+ bl[118] br[118] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_121 
+ bl[119] br[119] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_122 
+ bl[120] br[120] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_123 
+ bl[121] br[121] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_124 
+ bl[122] br[122] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_125 
+ bl[123] br[123] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_126 
+ bl[124] br[124] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_127 
+ bl[125] br[125] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_128 
+ bl[126] br[126] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_129 
+ bl[127] br[127] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_130 
+ vdd vdd vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_131 
+ vdd vdd vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_0 
+ vdd vdd vss vdd vpb vnb wl[31] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_33_1 
+ rbl rbr vss vdd vpb vnb wl[31] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_33_2 
+ bl[0] br[0] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_3 
+ bl[1] br[1] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_4 
+ bl[2] br[2] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_5 
+ bl[3] br[3] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_6 
+ bl[4] br[4] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_7 
+ bl[5] br[5] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_8 
+ bl[6] br[6] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_9 
+ bl[7] br[7] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_10 
+ bl[8] br[8] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_11 
+ bl[9] br[9] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_12 
+ bl[10] br[10] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_13 
+ bl[11] br[11] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_14 
+ bl[12] br[12] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_15 
+ bl[13] br[13] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_16 
+ bl[14] br[14] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_17 
+ bl[15] br[15] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_18 
+ bl[16] br[16] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_19 
+ bl[17] br[17] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_20 
+ bl[18] br[18] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_21 
+ bl[19] br[19] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_22 
+ bl[20] br[20] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_23 
+ bl[21] br[21] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_24 
+ bl[22] br[22] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_25 
+ bl[23] br[23] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_26 
+ bl[24] br[24] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_27 
+ bl[25] br[25] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_28 
+ bl[26] br[26] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_29 
+ bl[27] br[27] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_30 
+ bl[28] br[28] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_31 
+ bl[29] br[29] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_32 
+ bl[30] br[30] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_33 
+ bl[31] br[31] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_34 
+ bl[32] br[32] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_35 
+ bl[33] br[33] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_36 
+ bl[34] br[34] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_37 
+ bl[35] br[35] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_38 
+ bl[36] br[36] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_39 
+ bl[37] br[37] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_40 
+ bl[38] br[38] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_41 
+ bl[39] br[39] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_42 
+ bl[40] br[40] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_43 
+ bl[41] br[41] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_44 
+ bl[42] br[42] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_45 
+ bl[43] br[43] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_46 
+ bl[44] br[44] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_47 
+ bl[45] br[45] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_48 
+ bl[46] br[46] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_49 
+ bl[47] br[47] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_50 
+ bl[48] br[48] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_51 
+ bl[49] br[49] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_52 
+ bl[50] br[50] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_53 
+ bl[51] br[51] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_54 
+ bl[52] br[52] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_55 
+ bl[53] br[53] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_56 
+ bl[54] br[54] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_57 
+ bl[55] br[55] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_58 
+ bl[56] br[56] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_59 
+ bl[57] br[57] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_60 
+ bl[58] br[58] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_61 
+ bl[59] br[59] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_62 
+ bl[60] br[60] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_63 
+ bl[61] br[61] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_64 
+ bl[62] br[62] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_65 
+ bl[63] br[63] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_66 
+ bl[64] br[64] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_67 
+ bl[65] br[65] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_68 
+ bl[66] br[66] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_69 
+ bl[67] br[67] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_70 
+ bl[68] br[68] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_71 
+ bl[69] br[69] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_72 
+ bl[70] br[70] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_73 
+ bl[71] br[71] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_74 
+ bl[72] br[72] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_75 
+ bl[73] br[73] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_76 
+ bl[74] br[74] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_77 
+ bl[75] br[75] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_78 
+ bl[76] br[76] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_79 
+ bl[77] br[77] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_80 
+ bl[78] br[78] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_81 
+ bl[79] br[79] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_82 
+ bl[80] br[80] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_83 
+ bl[81] br[81] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_84 
+ bl[82] br[82] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_85 
+ bl[83] br[83] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_86 
+ bl[84] br[84] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_87 
+ bl[85] br[85] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_88 
+ bl[86] br[86] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_89 
+ bl[87] br[87] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_90 
+ bl[88] br[88] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_91 
+ bl[89] br[89] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_92 
+ bl[90] br[90] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_93 
+ bl[91] br[91] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_94 
+ bl[92] br[92] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_95 
+ bl[93] br[93] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_96 
+ bl[94] br[94] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_97 
+ bl[95] br[95] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_98 
+ bl[96] br[96] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_99 
+ bl[97] br[97] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_100 
+ bl[98] br[98] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_101 
+ bl[99] br[99] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_102 
+ bl[100] br[100] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_103 
+ bl[101] br[101] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_104 
+ bl[102] br[102] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_105 
+ bl[103] br[103] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_106 
+ bl[104] br[104] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_107 
+ bl[105] br[105] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_108 
+ bl[106] br[106] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_109 
+ bl[107] br[107] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_110 
+ bl[108] br[108] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_111 
+ bl[109] br[109] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_112 
+ bl[110] br[110] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_113 
+ bl[111] br[111] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_114 
+ bl[112] br[112] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_115 
+ bl[113] br[113] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_116 
+ bl[114] br[114] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_117 
+ bl[115] br[115] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_118 
+ bl[116] br[116] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_119 
+ bl[117] br[117] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_120 
+ bl[118] br[118] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_121 
+ bl[119] br[119] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_122 
+ bl[120] br[120] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_123 
+ bl[121] br[121] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_124 
+ bl[122] br[122] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_125 
+ bl[123] br[123] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_126 
+ bl[124] br[124] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_127 
+ bl[125] br[125] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_128 
+ bl[126] br[126] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_129 
+ bl[127] br[127] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_130 
+ vdd vdd vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_131 
+ vdd vdd vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_0 
+ vdd vdd vss vdd vpb vnb wl[32] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_34_1 
+ rbl rbr vss vdd vpb vnb wl[32] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_34_2 
+ bl[0] br[0] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_3 
+ bl[1] br[1] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_4 
+ bl[2] br[2] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_5 
+ bl[3] br[3] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_6 
+ bl[4] br[4] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_7 
+ bl[5] br[5] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_8 
+ bl[6] br[6] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_9 
+ bl[7] br[7] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_10 
+ bl[8] br[8] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_11 
+ bl[9] br[9] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_12 
+ bl[10] br[10] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_13 
+ bl[11] br[11] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_14 
+ bl[12] br[12] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_15 
+ bl[13] br[13] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_16 
+ bl[14] br[14] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_17 
+ bl[15] br[15] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_18 
+ bl[16] br[16] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_19 
+ bl[17] br[17] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_20 
+ bl[18] br[18] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_21 
+ bl[19] br[19] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_22 
+ bl[20] br[20] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_23 
+ bl[21] br[21] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_24 
+ bl[22] br[22] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_25 
+ bl[23] br[23] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_26 
+ bl[24] br[24] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_27 
+ bl[25] br[25] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_28 
+ bl[26] br[26] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_29 
+ bl[27] br[27] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_30 
+ bl[28] br[28] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_31 
+ bl[29] br[29] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_32 
+ bl[30] br[30] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_33 
+ bl[31] br[31] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_34 
+ bl[32] br[32] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_35 
+ bl[33] br[33] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_36 
+ bl[34] br[34] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_37 
+ bl[35] br[35] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_38 
+ bl[36] br[36] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_39 
+ bl[37] br[37] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_40 
+ bl[38] br[38] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_41 
+ bl[39] br[39] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_42 
+ bl[40] br[40] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_43 
+ bl[41] br[41] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_44 
+ bl[42] br[42] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_45 
+ bl[43] br[43] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_46 
+ bl[44] br[44] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_47 
+ bl[45] br[45] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_48 
+ bl[46] br[46] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_49 
+ bl[47] br[47] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_50 
+ bl[48] br[48] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_51 
+ bl[49] br[49] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_52 
+ bl[50] br[50] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_53 
+ bl[51] br[51] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_54 
+ bl[52] br[52] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_55 
+ bl[53] br[53] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_56 
+ bl[54] br[54] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_57 
+ bl[55] br[55] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_58 
+ bl[56] br[56] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_59 
+ bl[57] br[57] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_60 
+ bl[58] br[58] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_61 
+ bl[59] br[59] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_62 
+ bl[60] br[60] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_63 
+ bl[61] br[61] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_64 
+ bl[62] br[62] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_65 
+ bl[63] br[63] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_66 
+ bl[64] br[64] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_67 
+ bl[65] br[65] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_68 
+ bl[66] br[66] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_69 
+ bl[67] br[67] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_70 
+ bl[68] br[68] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_71 
+ bl[69] br[69] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_72 
+ bl[70] br[70] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_73 
+ bl[71] br[71] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_74 
+ bl[72] br[72] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_75 
+ bl[73] br[73] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_76 
+ bl[74] br[74] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_77 
+ bl[75] br[75] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_78 
+ bl[76] br[76] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_79 
+ bl[77] br[77] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_80 
+ bl[78] br[78] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_81 
+ bl[79] br[79] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_82 
+ bl[80] br[80] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_83 
+ bl[81] br[81] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_84 
+ bl[82] br[82] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_85 
+ bl[83] br[83] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_86 
+ bl[84] br[84] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_87 
+ bl[85] br[85] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_88 
+ bl[86] br[86] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_89 
+ bl[87] br[87] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_90 
+ bl[88] br[88] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_91 
+ bl[89] br[89] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_92 
+ bl[90] br[90] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_93 
+ bl[91] br[91] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_94 
+ bl[92] br[92] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_95 
+ bl[93] br[93] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_96 
+ bl[94] br[94] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_97 
+ bl[95] br[95] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_98 
+ bl[96] br[96] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_99 
+ bl[97] br[97] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_100 
+ bl[98] br[98] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_101 
+ bl[99] br[99] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_102 
+ bl[100] br[100] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_103 
+ bl[101] br[101] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_104 
+ bl[102] br[102] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_105 
+ bl[103] br[103] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_106 
+ bl[104] br[104] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_107 
+ bl[105] br[105] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_108 
+ bl[106] br[106] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_109 
+ bl[107] br[107] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_110 
+ bl[108] br[108] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_111 
+ bl[109] br[109] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_112 
+ bl[110] br[110] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_113 
+ bl[111] br[111] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_114 
+ bl[112] br[112] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_115 
+ bl[113] br[113] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_116 
+ bl[114] br[114] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_117 
+ bl[115] br[115] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_118 
+ bl[116] br[116] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_119 
+ bl[117] br[117] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_120 
+ bl[118] br[118] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_121 
+ bl[119] br[119] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_122 
+ bl[120] br[120] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_123 
+ bl[121] br[121] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_124 
+ bl[122] br[122] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_125 
+ bl[123] br[123] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_126 
+ bl[124] br[124] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_127 
+ bl[125] br[125] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_128 
+ bl[126] br[126] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_129 
+ bl[127] br[127] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_130 
+ vdd vdd vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_131 
+ vdd vdd vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_0 
+ vdd vdd vss vdd vpb vnb wl[33] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_35_1 
+ rbl rbr vss vdd vpb vnb wl[33] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_35_2 
+ bl[0] br[0] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_3 
+ bl[1] br[1] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_4 
+ bl[2] br[2] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_5 
+ bl[3] br[3] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_6 
+ bl[4] br[4] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_7 
+ bl[5] br[5] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_8 
+ bl[6] br[6] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_9 
+ bl[7] br[7] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_10 
+ bl[8] br[8] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_11 
+ bl[9] br[9] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_12 
+ bl[10] br[10] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_13 
+ bl[11] br[11] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_14 
+ bl[12] br[12] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_15 
+ bl[13] br[13] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_16 
+ bl[14] br[14] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_17 
+ bl[15] br[15] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_18 
+ bl[16] br[16] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_19 
+ bl[17] br[17] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_20 
+ bl[18] br[18] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_21 
+ bl[19] br[19] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_22 
+ bl[20] br[20] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_23 
+ bl[21] br[21] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_24 
+ bl[22] br[22] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_25 
+ bl[23] br[23] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_26 
+ bl[24] br[24] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_27 
+ bl[25] br[25] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_28 
+ bl[26] br[26] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_29 
+ bl[27] br[27] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_30 
+ bl[28] br[28] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_31 
+ bl[29] br[29] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_32 
+ bl[30] br[30] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_33 
+ bl[31] br[31] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_34 
+ bl[32] br[32] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_35 
+ bl[33] br[33] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_36 
+ bl[34] br[34] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_37 
+ bl[35] br[35] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_38 
+ bl[36] br[36] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_39 
+ bl[37] br[37] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_40 
+ bl[38] br[38] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_41 
+ bl[39] br[39] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_42 
+ bl[40] br[40] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_43 
+ bl[41] br[41] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_44 
+ bl[42] br[42] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_45 
+ bl[43] br[43] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_46 
+ bl[44] br[44] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_47 
+ bl[45] br[45] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_48 
+ bl[46] br[46] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_49 
+ bl[47] br[47] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_50 
+ bl[48] br[48] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_51 
+ bl[49] br[49] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_52 
+ bl[50] br[50] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_53 
+ bl[51] br[51] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_54 
+ bl[52] br[52] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_55 
+ bl[53] br[53] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_56 
+ bl[54] br[54] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_57 
+ bl[55] br[55] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_58 
+ bl[56] br[56] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_59 
+ bl[57] br[57] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_60 
+ bl[58] br[58] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_61 
+ bl[59] br[59] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_62 
+ bl[60] br[60] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_63 
+ bl[61] br[61] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_64 
+ bl[62] br[62] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_65 
+ bl[63] br[63] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_66 
+ bl[64] br[64] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_67 
+ bl[65] br[65] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_68 
+ bl[66] br[66] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_69 
+ bl[67] br[67] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_70 
+ bl[68] br[68] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_71 
+ bl[69] br[69] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_72 
+ bl[70] br[70] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_73 
+ bl[71] br[71] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_74 
+ bl[72] br[72] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_75 
+ bl[73] br[73] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_76 
+ bl[74] br[74] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_77 
+ bl[75] br[75] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_78 
+ bl[76] br[76] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_79 
+ bl[77] br[77] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_80 
+ bl[78] br[78] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_81 
+ bl[79] br[79] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_82 
+ bl[80] br[80] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_83 
+ bl[81] br[81] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_84 
+ bl[82] br[82] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_85 
+ bl[83] br[83] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_86 
+ bl[84] br[84] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_87 
+ bl[85] br[85] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_88 
+ bl[86] br[86] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_89 
+ bl[87] br[87] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_90 
+ bl[88] br[88] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_91 
+ bl[89] br[89] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_92 
+ bl[90] br[90] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_93 
+ bl[91] br[91] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_94 
+ bl[92] br[92] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_95 
+ bl[93] br[93] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_96 
+ bl[94] br[94] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_97 
+ bl[95] br[95] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_98 
+ bl[96] br[96] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_99 
+ bl[97] br[97] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_100 
+ bl[98] br[98] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_101 
+ bl[99] br[99] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_102 
+ bl[100] br[100] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_103 
+ bl[101] br[101] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_104 
+ bl[102] br[102] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_105 
+ bl[103] br[103] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_106 
+ bl[104] br[104] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_107 
+ bl[105] br[105] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_108 
+ bl[106] br[106] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_109 
+ bl[107] br[107] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_110 
+ bl[108] br[108] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_111 
+ bl[109] br[109] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_112 
+ bl[110] br[110] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_113 
+ bl[111] br[111] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_114 
+ bl[112] br[112] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_115 
+ bl[113] br[113] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_116 
+ bl[114] br[114] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_117 
+ bl[115] br[115] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_118 
+ bl[116] br[116] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_119 
+ bl[117] br[117] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_120 
+ bl[118] br[118] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_121 
+ bl[119] br[119] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_122 
+ bl[120] br[120] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_123 
+ bl[121] br[121] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_124 
+ bl[122] br[122] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_125 
+ bl[123] br[123] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_126 
+ bl[124] br[124] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_127 
+ bl[125] br[125] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_128 
+ bl[126] br[126] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_129 
+ bl[127] br[127] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_130 
+ vdd vdd vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_131 
+ vdd vdd vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_0 
+ vdd vdd vss vdd vpb vnb wl[34] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_36_1 
+ rbl rbr vss vdd vpb vnb wl[34] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_36_2 
+ bl[0] br[0] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_3 
+ bl[1] br[1] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_4 
+ bl[2] br[2] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_5 
+ bl[3] br[3] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_6 
+ bl[4] br[4] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_7 
+ bl[5] br[5] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_8 
+ bl[6] br[6] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_9 
+ bl[7] br[7] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_10 
+ bl[8] br[8] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_11 
+ bl[9] br[9] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_12 
+ bl[10] br[10] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_13 
+ bl[11] br[11] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_14 
+ bl[12] br[12] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_15 
+ bl[13] br[13] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_16 
+ bl[14] br[14] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_17 
+ bl[15] br[15] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_18 
+ bl[16] br[16] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_19 
+ bl[17] br[17] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_20 
+ bl[18] br[18] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_21 
+ bl[19] br[19] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_22 
+ bl[20] br[20] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_23 
+ bl[21] br[21] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_24 
+ bl[22] br[22] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_25 
+ bl[23] br[23] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_26 
+ bl[24] br[24] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_27 
+ bl[25] br[25] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_28 
+ bl[26] br[26] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_29 
+ bl[27] br[27] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_30 
+ bl[28] br[28] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_31 
+ bl[29] br[29] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_32 
+ bl[30] br[30] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_33 
+ bl[31] br[31] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_34 
+ bl[32] br[32] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_35 
+ bl[33] br[33] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_36 
+ bl[34] br[34] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_37 
+ bl[35] br[35] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_38 
+ bl[36] br[36] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_39 
+ bl[37] br[37] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_40 
+ bl[38] br[38] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_41 
+ bl[39] br[39] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_42 
+ bl[40] br[40] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_43 
+ bl[41] br[41] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_44 
+ bl[42] br[42] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_45 
+ bl[43] br[43] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_46 
+ bl[44] br[44] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_47 
+ bl[45] br[45] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_48 
+ bl[46] br[46] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_49 
+ bl[47] br[47] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_50 
+ bl[48] br[48] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_51 
+ bl[49] br[49] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_52 
+ bl[50] br[50] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_53 
+ bl[51] br[51] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_54 
+ bl[52] br[52] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_55 
+ bl[53] br[53] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_56 
+ bl[54] br[54] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_57 
+ bl[55] br[55] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_58 
+ bl[56] br[56] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_59 
+ bl[57] br[57] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_60 
+ bl[58] br[58] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_61 
+ bl[59] br[59] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_62 
+ bl[60] br[60] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_63 
+ bl[61] br[61] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_64 
+ bl[62] br[62] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_65 
+ bl[63] br[63] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_66 
+ bl[64] br[64] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_67 
+ bl[65] br[65] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_68 
+ bl[66] br[66] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_69 
+ bl[67] br[67] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_70 
+ bl[68] br[68] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_71 
+ bl[69] br[69] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_72 
+ bl[70] br[70] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_73 
+ bl[71] br[71] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_74 
+ bl[72] br[72] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_75 
+ bl[73] br[73] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_76 
+ bl[74] br[74] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_77 
+ bl[75] br[75] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_78 
+ bl[76] br[76] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_79 
+ bl[77] br[77] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_80 
+ bl[78] br[78] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_81 
+ bl[79] br[79] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_82 
+ bl[80] br[80] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_83 
+ bl[81] br[81] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_84 
+ bl[82] br[82] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_85 
+ bl[83] br[83] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_86 
+ bl[84] br[84] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_87 
+ bl[85] br[85] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_88 
+ bl[86] br[86] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_89 
+ bl[87] br[87] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_90 
+ bl[88] br[88] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_91 
+ bl[89] br[89] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_92 
+ bl[90] br[90] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_93 
+ bl[91] br[91] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_94 
+ bl[92] br[92] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_95 
+ bl[93] br[93] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_96 
+ bl[94] br[94] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_97 
+ bl[95] br[95] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_98 
+ bl[96] br[96] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_99 
+ bl[97] br[97] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_100 
+ bl[98] br[98] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_101 
+ bl[99] br[99] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_102 
+ bl[100] br[100] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_103 
+ bl[101] br[101] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_104 
+ bl[102] br[102] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_105 
+ bl[103] br[103] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_106 
+ bl[104] br[104] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_107 
+ bl[105] br[105] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_108 
+ bl[106] br[106] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_109 
+ bl[107] br[107] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_110 
+ bl[108] br[108] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_111 
+ bl[109] br[109] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_112 
+ bl[110] br[110] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_113 
+ bl[111] br[111] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_114 
+ bl[112] br[112] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_115 
+ bl[113] br[113] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_116 
+ bl[114] br[114] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_117 
+ bl[115] br[115] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_118 
+ bl[116] br[116] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_119 
+ bl[117] br[117] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_120 
+ bl[118] br[118] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_121 
+ bl[119] br[119] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_122 
+ bl[120] br[120] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_123 
+ bl[121] br[121] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_124 
+ bl[122] br[122] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_125 
+ bl[123] br[123] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_126 
+ bl[124] br[124] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_127 
+ bl[125] br[125] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_128 
+ bl[126] br[126] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_129 
+ bl[127] br[127] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_130 
+ vdd vdd vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_131 
+ vdd vdd vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_0 
+ vdd vdd vss vdd vpb vnb wl[35] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_37_1 
+ rbl rbr vss vdd vpb vnb wl[35] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_37_2 
+ bl[0] br[0] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_3 
+ bl[1] br[1] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_4 
+ bl[2] br[2] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_5 
+ bl[3] br[3] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_6 
+ bl[4] br[4] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_7 
+ bl[5] br[5] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_8 
+ bl[6] br[6] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_9 
+ bl[7] br[7] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_10 
+ bl[8] br[8] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_11 
+ bl[9] br[9] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_12 
+ bl[10] br[10] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_13 
+ bl[11] br[11] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_14 
+ bl[12] br[12] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_15 
+ bl[13] br[13] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_16 
+ bl[14] br[14] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_17 
+ bl[15] br[15] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_18 
+ bl[16] br[16] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_19 
+ bl[17] br[17] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_20 
+ bl[18] br[18] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_21 
+ bl[19] br[19] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_22 
+ bl[20] br[20] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_23 
+ bl[21] br[21] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_24 
+ bl[22] br[22] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_25 
+ bl[23] br[23] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_26 
+ bl[24] br[24] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_27 
+ bl[25] br[25] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_28 
+ bl[26] br[26] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_29 
+ bl[27] br[27] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_30 
+ bl[28] br[28] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_31 
+ bl[29] br[29] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_32 
+ bl[30] br[30] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_33 
+ bl[31] br[31] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_34 
+ bl[32] br[32] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_35 
+ bl[33] br[33] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_36 
+ bl[34] br[34] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_37 
+ bl[35] br[35] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_38 
+ bl[36] br[36] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_39 
+ bl[37] br[37] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_40 
+ bl[38] br[38] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_41 
+ bl[39] br[39] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_42 
+ bl[40] br[40] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_43 
+ bl[41] br[41] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_44 
+ bl[42] br[42] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_45 
+ bl[43] br[43] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_46 
+ bl[44] br[44] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_47 
+ bl[45] br[45] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_48 
+ bl[46] br[46] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_49 
+ bl[47] br[47] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_50 
+ bl[48] br[48] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_51 
+ bl[49] br[49] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_52 
+ bl[50] br[50] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_53 
+ bl[51] br[51] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_54 
+ bl[52] br[52] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_55 
+ bl[53] br[53] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_56 
+ bl[54] br[54] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_57 
+ bl[55] br[55] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_58 
+ bl[56] br[56] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_59 
+ bl[57] br[57] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_60 
+ bl[58] br[58] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_61 
+ bl[59] br[59] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_62 
+ bl[60] br[60] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_63 
+ bl[61] br[61] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_64 
+ bl[62] br[62] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_65 
+ bl[63] br[63] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_66 
+ bl[64] br[64] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_67 
+ bl[65] br[65] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_68 
+ bl[66] br[66] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_69 
+ bl[67] br[67] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_70 
+ bl[68] br[68] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_71 
+ bl[69] br[69] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_72 
+ bl[70] br[70] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_73 
+ bl[71] br[71] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_74 
+ bl[72] br[72] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_75 
+ bl[73] br[73] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_76 
+ bl[74] br[74] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_77 
+ bl[75] br[75] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_78 
+ bl[76] br[76] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_79 
+ bl[77] br[77] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_80 
+ bl[78] br[78] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_81 
+ bl[79] br[79] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_82 
+ bl[80] br[80] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_83 
+ bl[81] br[81] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_84 
+ bl[82] br[82] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_85 
+ bl[83] br[83] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_86 
+ bl[84] br[84] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_87 
+ bl[85] br[85] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_88 
+ bl[86] br[86] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_89 
+ bl[87] br[87] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_90 
+ bl[88] br[88] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_91 
+ bl[89] br[89] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_92 
+ bl[90] br[90] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_93 
+ bl[91] br[91] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_94 
+ bl[92] br[92] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_95 
+ bl[93] br[93] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_96 
+ bl[94] br[94] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_97 
+ bl[95] br[95] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_98 
+ bl[96] br[96] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_99 
+ bl[97] br[97] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_100 
+ bl[98] br[98] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_101 
+ bl[99] br[99] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_102 
+ bl[100] br[100] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_103 
+ bl[101] br[101] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_104 
+ bl[102] br[102] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_105 
+ bl[103] br[103] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_106 
+ bl[104] br[104] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_107 
+ bl[105] br[105] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_108 
+ bl[106] br[106] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_109 
+ bl[107] br[107] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_110 
+ bl[108] br[108] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_111 
+ bl[109] br[109] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_112 
+ bl[110] br[110] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_113 
+ bl[111] br[111] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_114 
+ bl[112] br[112] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_115 
+ bl[113] br[113] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_116 
+ bl[114] br[114] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_117 
+ bl[115] br[115] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_118 
+ bl[116] br[116] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_119 
+ bl[117] br[117] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_120 
+ bl[118] br[118] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_121 
+ bl[119] br[119] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_122 
+ bl[120] br[120] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_123 
+ bl[121] br[121] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_124 
+ bl[122] br[122] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_125 
+ bl[123] br[123] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_126 
+ bl[124] br[124] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_127 
+ bl[125] br[125] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_128 
+ bl[126] br[126] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_129 
+ bl[127] br[127] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_130 
+ vdd vdd vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_131 
+ vdd vdd vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_0 
+ vdd vdd vss vdd vpb vnb wl[36] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_38_1 
+ rbl rbr vss vdd vpb vnb wl[36] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_38_2 
+ bl[0] br[0] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_3 
+ bl[1] br[1] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_4 
+ bl[2] br[2] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_5 
+ bl[3] br[3] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_6 
+ bl[4] br[4] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_7 
+ bl[5] br[5] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_8 
+ bl[6] br[6] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_9 
+ bl[7] br[7] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_10 
+ bl[8] br[8] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_11 
+ bl[9] br[9] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_12 
+ bl[10] br[10] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_13 
+ bl[11] br[11] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_14 
+ bl[12] br[12] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_15 
+ bl[13] br[13] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_16 
+ bl[14] br[14] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_17 
+ bl[15] br[15] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_18 
+ bl[16] br[16] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_19 
+ bl[17] br[17] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_20 
+ bl[18] br[18] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_21 
+ bl[19] br[19] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_22 
+ bl[20] br[20] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_23 
+ bl[21] br[21] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_24 
+ bl[22] br[22] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_25 
+ bl[23] br[23] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_26 
+ bl[24] br[24] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_27 
+ bl[25] br[25] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_28 
+ bl[26] br[26] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_29 
+ bl[27] br[27] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_30 
+ bl[28] br[28] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_31 
+ bl[29] br[29] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_32 
+ bl[30] br[30] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_33 
+ bl[31] br[31] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_34 
+ bl[32] br[32] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_35 
+ bl[33] br[33] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_36 
+ bl[34] br[34] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_37 
+ bl[35] br[35] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_38 
+ bl[36] br[36] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_39 
+ bl[37] br[37] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_40 
+ bl[38] br[38] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_41 
+ bl[39] br[39] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_42 
+ bl[40] br[40] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_43 
+ bl[41] br[41] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_44 
+ bl[42] br[42] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_45 
+ bl[43] br[43] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_46 
+ bl[44] br[44] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_47 
+ bl[45] br[45] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_48 
+ bl[46] br[46] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_49 
+ bl[47] br[47] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_50 
+ bl[48] br[48] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_51 
+ bl[49] br[49] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_52 
+ bl[50] br[50] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_53 
+ bl[51] br[51] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_54 
+ bl[52] br[52] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_55 
+ bl[53] br[53] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_56 
+ bl[54] br[54] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_57 
+ bl[55] br[55] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_58 
+ bl[56] br[56] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_59 
+ bl[57] br[57] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_60 
+ bl[58] br[58] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_61 
+ bl[59] br[59] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_62 
+ bl[60] br[60] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_63 
+ bl[61] br[61] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_64 
+ bl[62] br[62] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_65 
+ bl[63] br[63] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_66 
+ bl[64] br[64] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_67 
+ bl[65] br[65] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_68 
+ bl[66] br[66] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_69 
+ bl[67] br[67] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_70 
+ bl[68] br[68] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_71 
+ bl[69] br[69] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_72 
+ bl[70] br[70] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_73 
+ bl[71] br[71] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_74 
+ bl[72] br[72] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_75 
+ bl[73] br[73] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_76 
+ bl[74] br[74] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_77 
+ bl[75] br[75] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_78 
+ bl[76] br[76] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_79 
+ bl[77] br[77] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_80 
+ bl[78] br[78] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_81 
+ bl[79] br[79] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_82 
+ bl[80] br[80] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_83 
+ bl[81] br[81] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_84 
+ bl[82] br[82] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_85 
+ bl[83] br[83] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_86 
+ bl[84] br[84] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_87 
+ bl[85] br[85] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_88 
+ bl[86] br[86] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_89 
+ bl[87] br[87] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_90 
+ bl[88] br[88] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_91 
+ bl[89] br[89] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_92 
+ bl[90] br[90] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_93 
+ bl[91] br[91] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_94 
+ bl[92] br[92] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_95 
+ bl[93] br[93] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_96 
+ bl[94] br[94] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_97 
+ bl[95] br[95] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_98 
+ bl[96] br[96] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_99 
+ bl[97] br[97] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_100 
+ bl[98] br[98] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_101 
+ bl[99] br[99] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_102 
+ bl[100] br[100] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_103 
+ bl[101] br[101] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_104 
+ bl[102] br[102] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_105 
+ bl[103] br[103] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_106 
+ bl[104] br[104] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_107 
+ bl[105] br[105] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_108 
+ bl[106] br[106] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_109 
+ bl[107] br[107] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_110 
+ bl[108] br[108] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_111 
+ bl[109] br[109] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_112 
+ bl[110] br[110] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_113 
+ bl[111] br[111] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_114 
+ bl[112] br[112] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_115 
+ bl[113] br[113] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_116 
+ bl[114] br[114] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_117 
+ bl[115] br[115] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_118 
+ bl[116] br[116] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_119 
+ bl[117] br[117] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_120 
+ bl[118] br[118] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_121 
+ bl[119] br[119] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_122 
+ bl[120] br[120] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_123 
+ bl[121] br[121] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_124 
+ bl[122] br[122] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_125 
+ bl[123] br[123] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_126 
+ bl[124] br[124] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_127 
+ bl[125] br[125] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_128 
+ bl[126] br[126] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_129 
+ bl[127] br[127] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_130 
+ vdd vdd vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_131 
+ vdd vdd vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_0 
+ vdd vdd vss vdd vpb vnb wl[37] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_39_1 
+ rbl rbr vss vdd vpb vnb wl[37] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_39_2 
+ bl[0] br[0] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_3 
+ bl[1] br[1] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_4 
+ bl[2] br[2] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_5 
+ bl[3] br[3] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_6 
+ bl[4] br[4] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_7 
+ bl[5] br[5] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_8 
+ bl[6] br[6] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_9 
+ bl[7] br[7] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_10 
+ bl[8] br[8] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_11 
+ bl[9] br[9] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_12 
+ bl[10] br[10] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_13 
+ bl[11] br[11] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_14 
+ bl[12] br[12] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_15 
+ bl[13] br[13] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_16 
+ bl[14] br[14] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_17 
+ bl[15] br[15] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_18 
+ bl[16] br[16] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_19 
+ bl[17] br[17] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_20 
+ bl[18] br[18] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_21 
+ bl[19] br[19] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_22 
+ bl[20] br[20] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_23 
+ bl[21] br[21] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_24 
+ bl[22] br[22] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_25 
+ bl[23] br[23] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_26 
+ bl[24] br[24] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_27 
+ bl[25] br[25] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_28 
+ bl[26] br[26] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_29 
+ bl[27] br[27] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_30 
+ bl[28] br[28] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_31 
+ bl[29] br[29] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_32 
+ bl[30] br[30] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_33 
+ bl[31] br[31] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_34 
+ bl[32] br[32] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_35 
+ bl[33] br[33] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_36 
+ bl[34] br[34] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_37 
+ bl[35] br[35] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_38 
+ bl[36] br[36] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_39 
+ bl[37] br[37] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_40 
+ bl[38] br[38] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_41 
+ bl[39] br[39] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_42 
+ bl[40] br[40] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_43 
+ bl[41] br[41] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_44 
+ bl[42] br[42] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_45 
+ bl[43] br[43] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_46 
+ bl[44] br[44] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_47 
+ bl[45] br[45] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_48 
+ bl[46] br[46] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_49 
+ bl[47] br[47] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_50 
+ bl[48] br[48] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_51 
+ bl[49] br[49] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_52 
+ bl[50] br[50] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_53 
+ bl[51] br[51] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_54 
+ bl[52] br[52] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_55 
+ bl[53] br[53] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_56 
+ bl[54] br[54] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_57 
+ bl[55] br[55] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_58 
+ bl[56] br[56] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_59 
+ bl[57] br[57] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_60 
+ bl[58] br[58] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_61 
+ bl[59] br[59] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_62 
+ bl[60] br[60] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_63 
+ bl[61] br[61] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_64 
+ bl[62] br[62] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_65 
+ bl[63] br[63] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_66 
+ bl[64] br[64] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_67 
+ bl[65] br[65] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_68 
+ bl[66] br[66] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_69 
+ bl[67] br[67] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_70 
+ bl[68] br[68] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_71 
+ bl[69] br[69] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_72 
+ bl[70] br[70] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_73 
+ bl[71] br[71] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_74 
+ bl[72] br[72] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_75 
+ bl[73] br[73] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_76 
+ bl[74] br[74] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_77 
+ bl[75] br[75] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_78 
+ bl[76] br[76] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_79 
+ bl[77] br[77] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_80 
+ bl[78] br[78] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_81 
+ bl[79] br[79] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_82 
+ bl[80] br[80] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_83 
+ bl[81] br[81] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_84 
+ bl[82] br[82] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_85 
+ bl[83] br[83] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_86 
+ bl[84] br[84] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_87 
+ bl[85] br[85] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_88 
+ bl[86] br[86] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_89 
+ bl[87] br[87] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_90 
+ bl[88] br[88] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_91 
+ bl[89] br[89] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_92 
+ bl[90] br[90] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_93 
+ bl[91] br[91] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_94 
+ bl[92] br[92] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_95 
+ bl[93] br[93] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_96 
+ bl[94] br[94] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_97 
+ bl[95] br[95] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_98 
+ bl[96] br[96] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_99 
+ bl[97] br[97] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_100 
+ bl[98] br[98] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_101 
+ bl[99] br[99] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_102 
+ bl[100] br[100] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_103 
+ bl[101] br[101] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_104 
+ bl[102] br[102] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_105 
+ bl[103] br[103] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_106 
+ bl[104] br[104] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_107 
+ bl[105] br[105] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_108 
+ bl[106] br[106] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_109 
+ bl[107] br[107] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_110 
+ bl[108] br[108] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_111 
+ bl[109] br[109] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_112 
+ bl[110] br[110] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_113 
+ bl[111] br[111] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_114 
+ bl[112] br[112] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_115 
+ bl[113] br[113] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_116 
+ bl[114] br[114] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_117 
+ bl[115] br[115] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_118 
+ bl[116] br[116] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_119 
+ bl[117] br[117] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_120 
+ bl[118] br[118] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_121 
+ bl[119] br[119] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_122 
+ bl[120] br[120] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_123 
+ bl[121] br[121] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_124 
+ bl[122] br[122] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_125 
+ bl[123] br[123] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_126 
+ bl[124] br[124] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_127 
+ bl[125] br[125] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_128 
+ bl[126] br[126] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_129 
+ bl[127] br[127] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_130 
+ vdd vdd vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_131 
+ vdd vdd vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_0 
+ vdd vdd vss vdd vpb vnb wl[38] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_40_1 
+ rbl rbr vss vdd vpb vnb wl[38] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_40_2 
+ bl[0] br[0] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_3 
+ bl[1] br[1] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_4 
+ bl[2] br[2] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_5 
+ bl[3] br[3] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_6 
+ bl[4] br[4] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_7 
+ bl[5] br[5] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_8 
+ bl[6] br[6] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_9 
+ bl[7] br[7] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_10 
+ bl[8] br[8] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_11 
+ bl[9] br[9] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_12 
+ bl[10] br[10] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_13 
+ bl[11] br[11] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_14 
+ bl[12] br[12] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_15 
+ bl[13] br[13] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_16 
+ bl[14] br[14] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_17 
+ bl[15] br[15] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_18 
+ bl[16] br[16] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_19 
+ bl[17] br[17] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_20 
+ bl[18] br[18] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_21 
+ bl[19] br[19] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_22 
+ bl[20] br[20] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_23 
+ bl[21] br[21] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_24 
+ bl[22] br[22] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_25 
+ bl[23] br[23] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_26 
+ bl[24] br[24] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_27 
+ bl[25] br[25] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_28 
+ bl[26] br[26] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_29 
+ bl[27] br[27] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_30 
+ bl[28] br[28] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_31 
+ bl[29] br[29] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_32 
+ bl[30] br[30] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_33 
+ bl[31] br[31] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_34 
+ bl[32] br[32] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_35 
+ bl[33] br[33] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_36 
+ bl[34] br[34] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_37 
+ bl[35] br[35] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_38 
+ bl[36] br[36] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_39 
+ bl[37] br[37] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_40 
+ bl[38] br[38] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_41 
+ bl[39] br[39] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_42 
+ bl[40] br[40] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_43 
+ bl[41] br[41] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_44 
+ bl[42] br[42] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_45 
+ bl[43] br[43] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_46 
+ bl[44] br[44] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_47 
+ bl[45] br[45] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_48 
+ bl[46] br[46] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_49 
+ bl[47] br[47] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_50 
+ bl[48] br[48] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_51 
+ bl[49] br[49] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_52 
+ bl[50] br[50] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_53 
+ bl[51] br[51] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_54 
+ bl[52] br[52] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_55 
+ bl[53] br[53] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_56 
+ bl[54] br[54] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_57 
+ bl[55] br[55] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_58 
+ bl[56] br[56] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_59 
+ bl[57] br[57] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_60 
+ bl[58] br[58] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_61 
+ bl[59] br[59] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_62 
+ bl[60] br[60] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_63 
+ bl[61] br[61] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_64 
+ bl[62] br[62] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_65 
+ bl[63] br[63] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_66 
+ bl[64] br[64] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_67 
+ bl[65] br[65] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_68 
+ bl[66] br[66] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_69 
+ bl[67] br[67] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_70 
+ bl[68] br[68] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_71 
+ bl[69] br[69] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_72 
+ bl[70] br[70] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_73 
+ bl[71] br[71] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_74 
+ bl[72] br[72] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_75 
+ bl[73] br[73] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_76 
+ bl[74] br[74] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_77 
+ bl[75] br[75] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_78 
+ bl[76] br[76] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_79 
+ bl[77] br[77] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_80 
+ bl[78] br[78] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_81 
+ bl[79] br[79] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_82 
+ bl[80] br[80] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_83 
+ bl[81] br[81] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_84 
+ bl[82] br[82] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_85 
+ bl[83] br[83] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_86 
+ bl[84] br[84] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_87 
+ bl[85] br[85] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_88 
+ bl[86] br[86] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_89 
+ bl[87] br[87] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_90 
+ bl[88] br[88] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_91 
+ bl[89] br[89] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_92 
+ bl[90] br[90] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_93 
+ bl[91] br[91] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_94 
+ bl[92] br[92] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_95 
+ bl[93] br[93] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_96 
+ bl[94] br[94] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_97 
+ bl[95] br[95] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_98 
+ bl[96] br[96] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_99 
+ bl[97] br[97] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_100 
+ bl[98] br[98] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_101 
+ bl[99] br[99] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_102 
+ bl[100] br[100] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_103 
+ bl[101] br[101] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_104 
+ bl[102] br[102] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_105 
+ bl[103] br[103] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_106 
+ bl[104] br[104] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_107 
+ bl[105] br[105] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_108 
+ bl[106] br[106] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_109 
+ bl[107] br[107] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_110 
+ bl[108] br[108] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_111 
+ bl[109] br[109] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_112 
+ bl[110] br[110] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_113 
+ bl[111] br[111] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_114 
+ bl[112] br[112] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_115 
+ bl[113] br[113] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_116 
+ bl[114] br[114] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_117 
+ bl[115] br[115] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_118 
+ bl[116] br[116] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_119 
+ bl[117] br[117] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_120 
+ bl[118] br[118] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_121 
+ bl[119] br[119] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_122 
+ bl[120] br[120] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_123 
+ bl[121] br[121] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_124 
+ bl[122] br[122] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_125 
+ bl[123] br[123] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_126 
+ bl[124] br[124] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_127 
+ bl[125] br[125] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_128 
+ bl[126] br[126] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_129 
+ bl[127] br[127] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_130 
+ vdd vdd vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_131 
+ vdd vdd vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_0 
+ vdd vdd vss vdd vpb vnb wl[39] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_41_1 
+ rbl rbr vss vdd vpb vnb wl[39] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_41_2 
+ bl[0] br[0] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_3 
+ bl[1] br[1] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_4 
+ bl[2] br[2] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_5 
+ bl[3] br[3] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_6 
+ bl[4] br[4] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_7 
+ bl[5] br[5] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_8 
+ bl[6] br[6] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_9 
+ bl[7] br[7] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_10 
+ bl[8] br[8] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_11 
+ bl[9] br[9] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_12 
+ bl[10] br[10] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_13 
+ bl[11] br[11] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_14 
+ bl[12] br[12] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_15 
+ bl[13] br[13] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_16 
+ bl[14] br[14] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_17 
+ bl[15] br[15] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_18 
+ bl[16] br[16] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_19 
+ bl[17] br[17] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_20 
+ bl[18] br[18] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_21 
+ bl[19] br[19] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_22 
+ bl[20] br[20] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_23 
+ bl[21] br[21] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_24 
+ bl[22] br[22] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_25 
+ bl[23] br[23] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_26 
+ bl[24] br[24] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_27 
+ bl[25] br[25] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_28 
+ bl[26] br[26] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_29 
+ bl[27] br[27] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_30 
+ bl[28] br[28] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_31 
+ bl[29] br[29] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_32 
+ bl[30] br[30] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_33 
+ bl[31] br[31] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_34 
+ bl[32] br[32] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_35 
+ bl[33] br[33] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_36 
+ bl[34] br[34] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_37 
+ bl[35] br[35] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_38 
+ bl[36] br[36] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_39 
+ bl[37] br[37] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_40 
+ bl[38] br[38] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_41 
+ bl[39] br[39] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_42 
+ bl[40] br[40] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_43 
+ bl[41] br[41] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_44 
+ bl[42] br[42] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_45 
+ bl[43] br[43] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_46 
+ bl[44] br[44] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_47 
+ bl[45] br[45] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_48 
+ bl[46] br[46] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_49 
+ bl[47] br[47] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_50 
+ bl[48] br[48] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_51 
+ bl[49] br[49] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_52 
+ bl[50] br[50] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_53 
+ bl[51] br[51] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_54 
+ bl[52] br[52] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_55 
+ bl[53] br[53] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_56 
+ bl[54] br[54] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_57 
+ bl[55] br[55] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_58 
+ bl[56] br[56] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_59 
+ bl[57] br[57] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_60 
+ bl[58] br[58] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_61 
+ bl[59] br[59] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_62 
+ bl[60] br[60] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_63 
+ bl[61] br[61] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_64 
+ bl[62] br[62] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_65 
+ bl[63] br[63] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_66 
+ bl[64] br[64] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_67 
+ bl[65] br[65] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_68 
+ bl[66] br[66] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_69 
+ bl[67] br[67] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_70 
+ bl[68] br[68] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_71 
+ bl[69] br[69] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_72 
+ bl[70] br[70] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_73 
+ bl[71] br[71] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_74 
+ bl[72] br[72] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_75 
+ bl[73] br[73] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_76 
+ bl[74] br[74] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_77 
+ bl[75] br[75] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_78 
+ bl[76] br[76] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_79 
+ bl[77] br[77] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_80 
+ bl[78] br[78] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_81 
+ bl[79] br[79] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_82 
+ bl[80] br[80] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_83 
+ bl[81] br[81] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_84 
+ bl[82] br[82] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_85 
+ bl[83] br[83] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_86 
+ bl[84] br[84] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_87 
+ bl[85] br[85] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_88 
+ bl[86] br[86] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_89 
+ bl[87] br[87] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_90 
+ bl[88] br[88] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_91 
+ bl[89] br[89] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_92 
+ bl[90] br[90] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_93 
+ bl[91] br[91] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_94 
+ bl[92] br[92] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_95 
+ bl[93] br[93] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_96 
+ bl[94] br[94] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_97 
+ bl[95] br[95] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_98 
+ bl[96] br[96] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_99 
+ bl[97] br[97] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_100 
+ bl[98] br[98] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_101 
+ bl[99] br[99] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_102 
+ bl[100] br[100] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_103 
+ bl[101] br[101] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_104 
+ bl[102] br[102] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_105 
+ bl[103] br[103] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_106 
+ bl[104] br[104] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_107 
+ bl[105] br[105] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_108 
+ bl[106] br[106] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_109 
+ bl[107] br[107] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_110 
+ bl[108] br[108] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_111 
+ bl[109] br[109] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_112 
+ bl[110] br[110] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_113 
+ bl[111] br[111] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_114 
+ bl[112] br[112] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_115 
+ bl[113] br[113] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_116 
+ bl[114] br[114] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_117 
+ bl[115] br[115] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_118 
+ bl[116] br[116] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_119 
+ bl[117] br[117] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_120 
+ bl[118] br[118] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_121 
+ bl[119] br[119] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_122 
+ bl[120] br[120] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_123 
+ bl[121] br[121] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_124 
+ bl[122] br[122] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_125 
+ bl[123] br[123] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_126 
+ bl[124] br[124] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_127 
+ bl[125] br[125] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_128 
+ bl[126] br[126] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_129 
+ bl[127] br[127] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_130 
+ vdd vdd vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_131 
+ vdd vdd vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_0 
+ vdd vdd vss vdd vpb vnb wl[40] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_42_1 
+ rbl rbr vss vdd vpb vnb wl[40] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_42_2 
+ bl[0] br[0] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_3 
+ bl[1] br[1] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_4 
+ bl[2] br[2] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_5 
+ bl[3] br[3] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_6 
+ bl[4] br[4] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_7 
+ bl[5] br[5] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_8 
+ bl[6] br[6] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_9 
+ bl[7] br[7] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_10 
+ bl[8] br[8] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_11 
+ bl[9] br[9] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_12 
+ bl[10] br[10] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_13 
+ bl[11] br[11] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_14 
+ bl[12] br[12] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_15 
+ bl[13] br[13] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_16 
+ bl[14] br[14] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_17 
+ bl[15] br[15] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_18 
+ bl[16] br[16] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_19 
+ bl[17] br[17] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_20 
+ bl[18] br[18] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_21 
+ bl[19] br[19] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_22 
+ bl[20] br[20] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_23 
+ bl[21] br[21] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_24 
+ bl[22] br[22] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_25 
+ bl[23] br[23] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_26 
+ bl[24] br[24] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_27 
+ bl[25] br[25] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_28 
+ bl[26] br[26] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_29 
+ bl[27] br[27] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_30 
+ bl[28] br[28] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_31 
+ bl[29] br[29] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_32 
+ bl[30] br[30] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_33 
+ bl[31] br[31] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_34 
+ bl[32] br[32] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_35 
+ bl[33] br[33] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_36 
+ bl[34] br[34] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_37 
+ bl[35] br[35] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_38 
+ bl[36] br[36] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_39 
+ bl[37] br[37] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_40 
+ bl[38] br[38] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_41 
+ bl[39] br[39] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_42 
+ bl[40] br[40] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_43 
+ bl[41] br[41] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_44 
+ bl[42] br[42] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_45 
+ bl[43] br[43] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_46 
+ bl[44] br[44] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_47 
+ bl[45] br[45] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_48 
+ bl[46] br[46] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_49 
+ bl[47] br[47] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_50 
+ bl[48] br[48] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_51 
+ bl[49] br[49] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_52 
+ bl[50] br[50] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_53 
+ bl[51] br[51] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_54 
+ bl[52] br[52] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_55 
+ bl[53] br[53] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_56 
+ bl[54] br[54] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_57 
+ bl[55] br[55] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_58 
+ bl[56] br[56] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_59 
+ bl[57] br[57] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_60 
+ bl[58] br[58] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_61 
+ bl[59] br[59] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_62 
+ bl[60] br[60] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_63 
+ bl[61] br[61] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_64 
+ bl[62] br[62] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_65 
+ bl[63] br[63] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_66 
+ bl[64] br[64] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_67 
+ bl[65] br[65] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_68 
+ bl[66] br[66] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_69 
+ bl[67] br[67] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_70 
+ bl[68] br[68] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_71 
+ bl[69] br[69] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_72 
+ bl[70] br[70] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_73 
+ bl[71] br[71] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_74 
+ bl[72] br[72] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_75 
+ bl[73] br[73] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_76 
+ bl[74] br[74] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_77 
+ bl[75] br[75] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_78 
+ bl[76] br[76] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_79 
+ bl[77] br[77] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_80 
+ bl[78] br[78] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_81 
+ bl[79] br[79] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_82 
+ bl[80] br[80] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_83 
+ bl[81] br[81] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_84 
+ bl[82] br[82] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_85 
+ bl[83] br[83] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_86 
+ bl[84] br[84] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_87 
+ bl[85] br[85] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_88 
+ bl[86] br[86] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_89 
+ bl[87] br[87] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_90 
+ bl[88] br[88] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_91 
+ bl[89] br[89] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_92 
+ bl[90] br[90] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_93 
+ bl[91] br[91] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_94 
+ bl[92] br[92] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_95 
+ bl[93] br[93] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_96 
+ bl[94] br[94] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_97 
+ bl[95] br[95] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_98 
+ bl[96] br[96] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_99 
+ bl[97] br[97] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_100 
+ bl[98] br[98] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_101 
+ bl[99] br[99] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_102 
+ bl[100] br[100] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_103 
+ bl[101] br[101] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_104 
+ bl[102] br[102] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_105 
+ bl[103] br[103] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_106 
+ bl[104] br[104] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_107 
+ bl[105] br[105] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_108 
+ bl[106] br[106] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_109 
+ bl[107] br[107] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_110 
+ bl[108] br[108] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_111 
+ bl[109] br[109] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_112 
+ bl[110] br[110] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_113 
+ bl[111] br[111] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_114 
+ bl[112] br[112] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_115 
+ bl[113] br[113] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_116 
+ bl[114] br[114] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_117 
+ bl[115] br[115] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_118 
+ bl[116] br[116] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_119 
+ bl[117] br[117] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_120 
+ bl[118] br[118] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_121 
+ bl[119] br[119] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_122 
+ bl[120] br[120] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_123 
+ bl[121] br[121] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_124 
+ bl[122] br[122] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_125 
+ bl[123] br[123] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_126 
+ bl[124] br[124] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_127 
+ bl[125] br[125] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_128 
+ bl[126] br[126] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_129 
+ bl[127] br[127] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_130 
+ vdd vdd vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_131 
+ vdd vdd vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_0 
+ vdd vdd vss vdd vpb vnb wl[41] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_43_1 
+ rbl rbr vss vdd vpb vnb wl[41] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_43_2 
+ bl[0] br[0] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_3 
+ bl[1] br[1] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_4 
+ bl[2] br[2] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_5 
+ bl[3] br[3] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_6 
+ bl[4] br[4] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_7 
+ bl[5] br[5] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_8 
+ bl[6] br[6] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_9 
+ bl[7] br[7] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_10 
+ bl[8] br[8] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_11 
+ bl[9] br[9] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_12 
+ bl[10] br[10] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_13 
+ bl[11] br[11] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_14 
+ bl[12] br[12] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_15 
+ bl[13] br[13] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_16 
+ bl[14] br[14] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_17 
+ bl[15] br[15] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_18 
+ bl[16] br[16] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_19 
+ bl[17] br[17] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_20 
+ bl[18] br[18] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_21 
+ bl[19] br[19] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_22 
+ bl[20] br[20] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_23 
+ bl[21] br[21] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_24 
+ bl[22] br[22] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_25 
+ bl[23] br[23] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_26 
+ bl[24] br[24] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_27 
+ bl[25] br[25] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_28 
+ bl[26] br[26] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_29 
+ bl[27] br[27] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_30 
+ bl[28] br[28] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_31 
+ bl[29] br[29] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_32 
+ bl[30] br[30] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_33 
+ bl[31] br[31] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_34 
+ bl[32] br[32] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_35 
+ bl[33] br[33] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_36 
+ bl[34] br[34] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_37 
+ bl[35] br[35] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_38 
+ bl[36] br[36] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_39 
+ bl[37] br[37] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_40 
+ bl[38] br[38] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_41 
+ bl[39] br[39] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_42 
+ bl[40] br[40] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_43 
+ bl[41] br[41] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_44 
+ bl[42] br[42] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_45 
+ bl[43] br[43] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_46 
+ bl[44] br[44] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_47 
+ bl[45] br[45] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_48 
+ bl[46] br[46] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_49 
+ bl[47] br[47] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_50 
+ bl[48] br[48] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_51 
+ bl[49] br[49] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_52 
+ bl[50] br[50] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_53 
+ bl[51] br[51] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_54 
+ bl[52] br[52] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_55 
+ bl[53] br[53] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_56 
+ bl[54] br[54] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_57 
+ bl[55] br[55] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_58 
+ bl[56] br[56] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_59 
+ bl[57] br[57] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_60 
+ bl[58] br[58] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_61 
+ bl[59] br[59] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_62 
+ bl[60] br[60] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_63 
+ bl[61] br[61] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_64 
+ bl[62] br[62] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_65 
+ bl[63] br[63] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_66 
+ bl[64] br[64] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_67 
+ bl[65] br[65] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_68 
+ bl[66] br[66] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_69 
+ bl[67] br[67] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_70 
+ bl[68] br[68] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_71 
+ bl[69] br[69] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_72 
+ bl[70] br[70] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_73 
+ bl[71] br[71] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_74 
+ bl[72] br[72] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_75 
+ bl[73] br[73] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_76 
+ bl[74] br[74] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_77 
+ bl[75] br[75] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_78 
+ bl[76] br[76] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_79 
+ bl[77] br[77] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_80 
+ bl[78] br[78] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_81 
+ bl[79] br[79] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_82 
+ bl[80] br[80] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_83 
+ bl[81] br[81] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_84 
+ bl[82] br[82] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_85 
+ bl[83] br[83] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_86 
+ bl[84] br[84] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_87 
+ bl[85] br[85] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_88 
+ bl[86] br[86] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_89 
+ bl[87] br[87] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_90 
+ bl[88] br[88] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_91 
+ bl[89] br[89] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_92 
+ bl[90] br[90] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_93 
+ bl[91] br[91] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_94 
+ bl[92] br[92] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_95 
+ bl[93] br[93] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_96 
+ bl[94] br[94] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_97 
+ bl[95] br[95] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_98 
+ bl[96] br[96] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_99 
+ bl[97] br[97] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_100 
+ bl[98] br[98] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_101 
+ bl[99] br[99] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_102 
+ bl[100] br[100] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_103 
+ bl[101] br[101] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_104 
+ bl[102] br[102] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_105 
+ bl[103] br[103] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_106 
+ bl[104] br[104] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_107 
+ bl[105] br[105] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_108 
+ bl[106] br[106] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_109 
+ bl[107] br[107] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_110 
+ bl[108] br[108] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_111 
+ bl[109] br[109] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_112 
+ bl[110] br[110] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_113 
+ bl[111] br[111] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_114 
+ bl[112] br[112] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_115 
+ bl[113] br[113] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_116 
+ bl[114] br[114] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_117 
+ bl[115] br[115] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_118 
+ bl[116] br[116] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_119 
+ bl[117] br[117] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_120 
+ bl[118] br[118] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_121 
+ bl[119] br[119] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_122 
+ bl[120] br[120] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_123 
+ bl[121] br[121] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_124 
+ bl[122] br[122] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_125 
+ bl[123] br[123] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_126 
+ bl[124] br[124] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_127 
+ bl[125] br[125] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_128 
+ bl[126] br[126] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_129 
+ bl[127] br[127] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_130 
+ vdd vdd vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_131 
+ vdd vdd vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_0 
+ vdd vdd vss vdd vpb vnb wl[42] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_44_1 
+ rbl rbr vss vdd vpb vnb wl[42] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_44_2 
+ bl[0] br[0] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_3 
+ bl[1] br[1] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_4 
+ bl[2] br[2] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_5 
+ bl[3] br[3] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_6 
+ bl[4] br[4] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_7 
+ bl[5] br[5] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_8 
+ bl[6] br[6] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_9 
+ bl[7] br[7] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_10 
+ bl[8] br[8] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_11 
+ bl[9] br[9] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_12 
+ bl[10] br[10] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_13 
+ bl[11] br[11] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_14 
+ bl[12] br[12] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_15 
+ bl[13] br[13] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_16 
+ bl[14] br[14] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_17 
+ bl[15] br[15] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_18 
+ bl[16] br[16] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_19 
+ bl[17] br[17] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_20 
+ bl[18] br[18] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_21 
+ bl[19] br[19] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_22 
+ bl[20] br[20] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_23 
+ bl[21] br[21] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_24 
+ bl[22] br[22] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_25 
+ bl[23] br[23] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_26 
+ bl[24] br[24] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_27 
+ bl[25] br[25] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_28 
+ bl[26] br[26] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_29 
+ bl[27] br[27] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_30 
+ bl[28] br[28] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_31 
+ bl[29] br[29] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_32 
+ bl[30] br[30] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_33 
+ bl[31] br[31] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_34 
+ bl[32] br[32] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_35 
+ bl[33] br[33] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_36 
+ bl[34] br[34] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_37 
+ bl[35] br[35] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_38 
+ bl[36] br[36] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_39 
+ bl[37] br[37] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_40 
+ bl[38] br[38] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_41 
+ bl[39] br[39] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_42 
+ bl[40] br[40] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_43 
+ bl[41] br[41] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_44 
+ bl[42] br[42] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_45 
+ bl[43] br[43] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_46 
+ bl[44] br[44] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_47 
+ bl[45] br[45] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_48 
+ bl[46] br[46] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_49 
+ bl[47] br[47] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_50 
+ bl[48] br[48] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_51 
+ bl[49] br[49] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_52 
+ bl[50] br[50] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_53 
+ bl[51] br[51] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_54 
+ bl[52] br[52] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_55 
+ bl[53] br[53] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_56 
+ bl[54] br[54] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_57 
+ bl[55] br[55] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_58 
+ bl[56] br[56] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_59 
+ bl[57] br[57] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_60 
+ bl[58] br[58] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_61 
+ bl[59] br[59] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_62 
+ bl[60] br[60] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_63 
+ bl[61] br[61] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_64 
+ bl[62] br[62] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_65 
+ bl[63] br[63] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_66 
+ bl[64] br[64] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_67 
+ bl[65] br[65] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_68 
+ bl[66] br[66] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_69 
+ bl[67] br[67] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_70 
+ bl[68] br[68] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_71 
+ bl[69] br[69] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_72 
+ bl[70] br[70] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_73 
+ bl[71] br[71] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_74 
+ bl[72] br[72] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_75 
+ bl[73] br[73] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_76 
+ bl[74] br[74] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_77 
+ bl[75] br[75] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_78 
+ bl[76] br[76] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_79 
+ bl[77] br[77] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_80 
+ bl[78] br[78] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_81 
+ bl[79] br[79] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_82 
+ bl[80] br[80] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_83 
+ bl[81] br[81] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_84 
+ bl[82] br[82] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_85 
+ bl[83] br[83] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_86 
+ bl[84] br[84] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_87 
+ bl[85] br[85] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_88 
+ bl[86] br[86] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_89 
+ bl[87] br[87] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_90 
+ bl[88] br[88] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_91 
+ bl[89] br[89] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_92 
+ bl[90] br[90] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_93 
+ bl[91] br[91] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_94 
+ bl[92] br[92] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_95 
+ bl[93] br[93] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_96 
+ bl[94] br[94] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_97 
+ bl[95] br[95] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_98 
+ bl[96] br[96] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_99 
+ bl[97] br[97] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_100 
+ bl[98] br[98] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_101 
+ bl[99] br[99] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_102 
+ bl[100] br[100] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_103 
+ bl[101] br[101] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_104 
+ bl[102] br[102] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_105 
+ bl[103] br[103] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_106 
+ bl[104] br[104] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_107 
+ bl[105] br[105] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_108 
+ bl[106] br[106] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_109 
+ bl[107] br[107] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_110 
+ bl[108] br[108] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_111 
+ bl[109] br[109] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_112 
+ bl[110] br[110] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_113 
+ bl[111] br[111] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_114 
+ bl[112] br[112] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_115 
+ bl[113] br[113] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_116 
+ bl[114] br[114] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_117 
+ bl[115] br[115] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_118 
+ bl[116] br[116] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_119 
+ bl[117] br[117] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_120 
+ bl[118] br[118] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_121 
+ bl[119] br[119] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_122 
+ bl[120] br[120] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_123 
+ bl[121] br[121] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_124 
+ bl[122] br[122] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_125 
+ bl[123] br[123] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_126 
+ bl[124] br[124] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_127 
+ bl[125] br[125] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_128 
+ bl[126] br[126] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_129 
+ bl[127] br[127] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_130 
+ vdd vdd vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_131 
+ vdd vdd vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_0 
+ vdd vdd vss vdd vpb vnb wl[43] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_45_1 
+ rbl rbr vss vdd vpb vnb wl[43] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_45_2 
+ bl[0] br[0] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_3 
+ bl[1] br[1] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_4 
+ bl[2] br[2] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_5 
+ bl[3] br[3] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_6 
+ bl[4] br[4] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_7 
+ bl[5] br[5] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_8 
+ bl[6] br[6] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_9 
+ bl[7] br[7] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_10 
+ bl[8] br[8] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_11 
+ bl[9] br[9] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_12 
+ bl[10] br[10] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_13 
+ bl[11] br[11] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_14 
+ bl[12] br[12] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_15 
+ bl[13] br[13] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_16 
+ bl[14] br[14] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_17 
+ bl[15] br[15] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_18 
+ bl[16] br[16] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_19 
+ bl[17] br[17] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_20 
+ bl[18] br[18] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_21 
+ bl[19] br[19] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_22 
+ bl[20] br[20] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_23 
+ bl[21] br[21] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_24 
+ bl[22] br[22] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_25 
+ bl[23] br[23] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_26 
+ bl[24] br[24] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_27 
+ bl[25] br[25] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_28 
+ bl[26] br[26] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_29 
+ bl[27] br[27] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_30 
+ bl[28] br[28] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_31 
+ bl[29] br[29] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_32 
+ bl[30] br[30] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_33 
+ bl[31] br[31] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_34 
+ bl[32] br[32] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_35 
+ bl[33] br[33] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_36 
+ bl[34] br[34] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_37 
+ bl[35] br[35] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_38 
+ bl[36] br[36] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_39 
+ bl[37] br[37] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_40 
+ bl[38] br[38] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_41 
+ bl[39] br[39] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_42 
+ bl[40] br[40] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_43 
+ bl[41] br[41] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_44 
+ bl[42] br[42] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_45 
+ bl[43] br[43] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_46 
+ bl[44] br[44] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_47 
+ bl[45] br[45] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_48 
+ bl[46] br[46] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_49 
+ bl[47] br[47] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_50 
+ bl[48] br[48] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_51 
+ bl[49] br[49] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_52 
+ bl[50] br[50] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_53 
+ bl[51] br[51] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_54 
+ bl[52] br[52] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_55 
+ bl[53] br[53] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_56 
+ bl[54] br[54] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_57 
+ bl[55] br[55] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_58 
+ bl[56] br[56] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_59 
+ bl[57] br[57] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_60 
+ bl[58] br[58] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_61 
+ bl[59] br[59] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_62 
+ bl[60] br[60] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_63 
+ bl[61] br[61] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_64 
+ bl[62] br[62] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_65 
+ bl[63] br[63] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_66 
+ bl[64] br[64] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_67 
+ bl[65] br[65] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_68 
+ bl[66] br[66] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_69 
+ bl[67] br[67] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_70 
+ bl[68] br[68] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_71 
+ bl[69] br[69] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_72 
+ bl[70] br[70] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_73 
+ bl[71] br[71] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_74 
+ bl[72] br[72] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_75 
+ bl[73] br[73] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_76 
+ bl[74] br[74] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_77 
+ bl[75] br[75] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_78 
+ bl[76] br[76] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_79 
+ bl[77] br[77] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_80 
+ bl[78] br[78] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_81 
+ bl[79] br[79] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_82 
+ bl[80] br[80] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_83 
+ bl[81] br[81] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_84 
+ bl[82] br[82] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_85 
+ bl[83] br[83] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_86 
+ bl[84] br[84] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_87 
+ bl[85] br[85] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_88 
+ bl[86] br[86] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_89 
+ bl[87] br[87] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_90 
+ bl[88] br[88] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_91 
+ bl[89] br[89] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_92 
+ bl[90] br[90] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_93 
+ bl[91] br[91] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_94 
+ bl[92] br[92] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_95 
+ bl[93] br[93] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_96 
+ bl[94] br[94] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_97 
+ bl[95] br[95] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_98 
+ bl[96] br[96] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_99 
+ bl[97] br[97] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_100 
+ bl[98] br[98] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_101 
+ bl[99] br[99] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_102 
+ bl[100] br[100] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_103 
+ bl[101] br[101] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_104 
+ bl[102] br[102] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_105 
+ bl[103] br[103] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_106 
+ bl[104] br[104] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_107 
+ bl[105] br[105] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_108 
+ bl[106] br[106] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_109 
+ bl[107] br[107] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_110 
+ bl[108] br[108] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_111 
+ bl[109] br[109] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_112 
+ bl[110] br[110] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_113 
+ bl[111] br[111] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_114 
+ bl[112] br[112] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_115 
+ bl[113] br[113] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_116 
+ bl[114] br[114] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_117 
+ bl[115] br[115] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_118 
+ bl[116] br[116] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_119 
+ bl[117] br[117] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_120 
+ bl[118] br[118] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_121 
+ bl[119] br[119] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_122 
+ bl[120] br[120] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_123 
+ bl[121] br[121] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_124 
+ bl[122] br[122] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_125 
+ bl[123] br[123] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_126 
+ bl[124] br[124] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_127 
+ bl[125] br[125] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_128 
+ bl[126] br[126] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_129 
+ bl[127] br[127] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_130 
+ vdd vdd vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_131 
+ vdd vdd vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_0 
+ vdd vdd vss vdd vpb vnb wl[44] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_46_1 
+ rbl rbr vss vdd vpb vnb wl[44] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_46_2 
+ bl[0] br[0] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_3 
+ bl[1] br[1] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_4 
+ bl[2] br[2] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_5 
+ bl[3] br[3] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_6 
+ bl[4] br[4] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_7 
+ bl[5] br[5] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_8 
+ bl[6] br[6] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_9 
+ bl[7] br[7] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_10 
+ bl[8] br[8] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_11 
+ bl[9] br[9] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_12 
+ bl[10] br[10] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_13 
+ bl[11] br[11] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_14 
+ bl[12] br[12] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_15 
+ bl[13] br[13] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_16 
+ bl[14] br[14] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_17 
+ bl[15] br[15] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_18 
+ bl[16] br[16] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_19 
+ bl[17] br[17] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_20 
+ bl[18] br[18] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_21 
+ bl[19] br[19] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_22 
+ bl[20] br[20] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_23 
+ bl[21] br[21] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_24 
+ bl[22] br[22] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_25 
+ bl[23] br[23] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_26 
+ bl[24] br[24] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_27 
+ bl[25] br[25] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_28 
+ bl[26] br[26] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_29 
+ bl[27] br[27] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_30 
+ bl[28] br[28] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_31 
+ bl[29] br[29] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_32 
+ bl[30] br[30] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_33 
+ bl[31] br[31] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_34 
+ bl[32] br[32] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_35 
+ bl[33] br[33] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_36 
+ bl[34] br[34] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_37 
+ bl[35] br[35] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_38 
+ bl[36] br[36] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_39 
+ bl[37] br[37] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_40 
+ bl[38] br[38] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_41 
+ bl[39] br[39] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_42 
+ bl[40] br[40] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_43 
+ bl[41] br[41] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_44 
+ bl[42] br[42] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_45 
+ bl[43] br[43] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_46 
+ bl[44] br[44] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_47 
+ bl[45] br[45] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_48 
+ bl[46] br[46] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_49 
+ bl[47] br[47] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_50 
+ bl[48] br[48] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_51 
+ bl[49] br[49] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_52 
+ bl[50] br[50] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_53 
+ bl[51] br[51] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_54 
+ bl[52] br[52] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_55 
+ bl[53] br[53] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_56 
+ bl[54] br[54] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_57 
+ bl[55] br[55] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_58 
+ bl[56] br[56] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_59 
+ bl[57] br[57] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_60 
+ bl[58] br[58] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_61 
+ bl[59] br[59] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_62 
+ bl[60] br[60] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_63 
+ bl[61] br[61] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_64 
+ bl[62] br[62] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_65 
+ bl[63] br[63] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_66 
+ bl[64] br[64] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_67 
+ bl[65] br[65] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_68 
+ bl[66] br[66] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_69 
+ bl[67] br[67] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_70 
+ bl[68] br[68] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_71 
+ bl[69] br[69] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_72 
+ bl[70] br[70] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_73 
+ bl[71] br[71] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_74 
+ bl[72] br[72] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_75 
+ bl[73] br[73] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_76 
+ bl[74] br[74] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_77 
+ bl[75] br[75] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_78 
+ bl[76] br[76] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_79 
+ bl[77] br[77] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_80 
+ bl[78] br[78] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_81 
+ bl[79] br[79] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_82 
+ bl[80] br[80] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_83 
+ bl[81] br[81] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_84 
+ bl[82] br[82] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_85 
+ bl[83] br[83] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_86 
+ bl[84] br[84] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_87 
+ bl[85] br[85] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_88 
+ bl[86] br[86] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_89 
+ bl[87] br[87] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_90 
+ bl[88] br[88] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_91 
+ bl[89] br[89] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_92 
+ bl[90] br[90] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_93 
+ bl[91] br[91] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_94 
+ bl[92] br[92] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_95 
+ bl[93] br[93] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_96 
+ bl[94] br[94] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_97 
+ bl[95] br[95] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_98 
+ bl[96] br[96] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_99 
+ bl[97] br[97] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_100 
+ bl[98] br[98] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_101 
+ bl[99] br[99] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_102 
+ bl[100] br[100] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_103 
+ bl[101] br[101] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_104 
+ bl[102] br[102] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_105 
+ bl[103] br[103] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_106 
+ bl[104] br[104] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_107 
+ bl[105] br[105] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_108 
+ bl[106] br[106] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_109 
+ bl[107] br[107] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_110 
+ bl[108] br[108] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_111 
+ bl[109] br[109] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_112 
+ bl[110] br[110] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_113 
+ bl[111] br[111] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_114 
+ bl[112] br[112] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_115 
+ bl[113] br[113] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_116 
+ bl[114] br[114] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_117 
+ bl[115] br[115] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_118 
+ bl[116] br[116] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_119 
+ bl[117] br[117] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_120 
+ bl[118] br[118] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_121 
+ bl[119] br[119] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_122 
+ bl[120] br[120] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_123 
+ bl[121] br[121] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_124 
+ bl[122] br[122] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_125 
+ bl[123] br[123] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_126 
+ bl[124] br[124] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_127 
+ bl[125] br[125] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_128 
+ bl[126] br[126] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_129 
+ bl[127] br[127] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_130 
+ vdd vdd vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_131 
+ vdd vdd vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_0 
+ vdd vdd vss vdd vpb vnb wl[45] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_47_1 
+ rbl rbr vss vdd vpb vnb wl[45] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_47_2 
+ bl[0] br[0] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_3 
+ bl[1] br[1] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_4 
+ bl[2] br[2] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_5 
+ bl[3] br[3] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_6 
+ bl[4] br[4] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_7 
+ bl[5] br[5] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_8 
+ bl[6] br[6] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_9 
+ bl[7] br[7] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_10 
+ bl[8] br[8] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_11 
+ bl[9] br[9] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_12 
+ bl[10] br[10] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_13 
+ bl[11] br[11] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_14 
+ bl[12] br[12] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_15 
+ bl[13] br[13] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_16 
+ bl[14] br[14] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_17 
+ bl[15] br[15] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_18 
+ bl[16] br[16] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_19 
+ bl[17] br[17] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_20 
+ bl[18] br[18] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_21 
+ bl[19] br[19] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_22 
+ bl[20] br[20] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_23 
+ bl[21] br[21] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_24 
+ bl[22] br[22] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_25 
+ bl[23] br[23] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_26 
+ bl[24] br[24] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_27 
+ bl[25] br[25] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_28 
+ bl[26] br[26] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_29 
+ bl[27] br[27] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_30 
+ bl[28] br[28] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_31 
+ bl[29] br[29] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_32 
+ bl[30] br[30] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_33 
+ bl[31] br[31] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_34 
+ bl[32] br[32] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_35 
+ bl[33] br[33] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_36 
+ bl[34] br[34] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_37 
+ bl[35] br[35] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_38 
+ bl[36] br[36] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_39 
+ bl[37] br[37] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_40 
+ bl[38] br[38] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_41 
+ bl[39] br[39] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_42 
+ bl[40] br[40] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_43 
+ bl[41] br[41] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_44 
+ bl[42] br[42] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_45 
+ bl[43] br[43] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_46 
+ bl[44] br[44] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_47 
+ bl[45] br[45] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_48 
+ bl[46] br[46] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_49 
+ bl[47] br[47] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_50 
+ bl[48] br[48] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_51 
+ bl[49] br[49] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_52 
+ bl[50] br[50] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_53 
+ bl[51] br[51] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_54 
+ bl[52] br[52] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_55 
+ bl[53] br[53] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_56 
+ bl[54] br[54] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_57 
+ bl[55] br[55] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_58 
+ bl[56] br[56] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_59 
+ bl[57] br[57] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_60 
+ bl[58] br[58] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_61 
+ bl[59] br[59] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_62 
+ bl[60] br[60] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_63 
+ bl[61] br[61] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_64 
+ bl[62] br[62] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_65 
+ bl[63] br[63] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_66 
+ bl[64] br[64] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_67 
+ bl[65] br[65] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_68 
+ bl[66] br[66] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_69 
+ bl[67] br[67] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_70 
+ bl[68] br[68] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_71 
+ bl[69] br[69] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_72 
+ bl[70] br[70] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_73 
+ bl[71] br[71] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_74 
+ bl[72] br[72] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_75 
+ bl[73] br[73] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_76 
+ bl[74] br[74] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_77 
+ bl[75] br[75] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_78 
+ bl[76] br[76] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_79 
+ bl[77] br[77] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_80 
+ bl[78] br[78] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_81 
+ bl[79] br[79] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_82 
+ bl[80] br[80] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_83 
+ bl[81] br[81] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_84 
+ bl[82] br[82] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_85 
+ bl[83] br[83] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_86 
+ bl[84] br[84] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_87 
+ bl[85] br[85] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_88 
+ bl[86] br[86] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_89 
+ bl[87] br[87] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_90 
+ bl[88] br[88] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_91 
+ bl[89] br[89] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_92 
+ bl[90] br[90] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_93 
+ bl[91] br[91] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_94 
+ bl[92] br[92] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_95 
+ bl[93] br[93] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_96 
+ bl[94] br[94] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_97 
+ bl[95] br[95] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_98 
+ bl[96] br[96] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_99 
+ bl[97] br[97] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_100 
+ bl[98] br[98] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_101 
+ bl[99] br[99] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_102 
+ bl[100] br[100] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_103 
+ bl[101] br[101] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_104 
+ bl[102] br[102] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_105 
+ bl[103] br[103] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_106 
+ bl[104] br[104] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_107 
+ bl[105] br[105] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_108 
+ bl[106] br[106] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_109 
+ bl[107] br[107] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_110 
+ bl[108] br[108] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_111 
+ bl[109] br[109] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_112 
+ bl[110] br[110] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_113 
+ bl[111] br[111] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_114 
+ bl[112] br[112] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_115 
+ bl[113] br[113] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_116 
+ bl[114] br[114] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_117 
+ bl[115] br[115] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_118 
+ bl[116] br[116] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_119 
+ bl[117] br[117] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_120 
+ bl[118] br[118] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_121 
+ bl[119] br[119] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_122 
+ bl[120] br[120] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_123 
+ bl[121] br[121] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_124 
+ bl[122] br[122] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_125 
+ bl[123] br[123] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_126 
+ bl[124] br[124] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_127 
+ bl[125] br[125] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_128 
+ bl[126] br[126] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_129 
+ bl[127] br[127] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_130 
+ vdd vdd vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_131 
+ vdd vdd vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_0 
+ vdd vdd vss vdd vpb vnb wl[46] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_48_1 
+ rbl rbr vss vdd vpb vnb wl[46] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_48_2 
+ bl[0] br[0] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_3 
+ bl[1] br[1] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_4 
+ bl[2] br[2] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_5 
+ bl[3] br[3] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_6 
+ bl[4] br[4] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_7 
+ bl[5] br[5] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_8 
+ bl[6] br[6] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_9 
+ bl[7] br[7] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_10 
+ bl[8] br[8] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_11 
+ bl[9] br[9] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_12 
+ bl[10] br[10] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_13 
+ bl[11] br[11] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_14 
+ bl[12] br[12] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_15 
+ bl[13] br[13] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_16 
+ bl[14] br[14] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_17 
+ bl[15] br[15] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_18 
+ bl[16] br[16] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_19 
+ bl[17] br[17] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_20 
+ bl[18] br[18] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_21 
+ bl[19] br[19] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_22 
+ bl[20] br[20] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_23 
+ bl[21] br[21] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_24 
+ bl[22] br[22] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_25 
+ bl[23] br[23] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_26 
+ bl[24] br[24] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_27 
+ bl[25] br[25] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_28 
+ bl[26] br[26] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_29 
+ bl[27] br[27] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_30 
+ bl[28] br[28] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_31 
+ bl[29] br[29] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_32 
+ bl[30] br[30] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_33 
+ bl[31] br[31] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_34 
+ bl[32] br[32] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_35 
+ bl[33] br[33] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_36 
+ bl[34] br[34] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_37 
+ bl[35] br[35] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_38 
+ bl[36] br[36] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_39 
+ bl[37] br[37] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_40 
+ bl[38] br[38] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_41 
+ bl[39] br[39] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_42 
+ bl[40] br[40] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_43 
+ bl[41] br[41] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_44 
+ bl[42] br[42] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_45 
+ bl[43] br[43] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_46 
+ bl[44] br[44] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_47 
+ bl[45] br[45] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_48 
+ bl[46] br[46] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_49 
+ bl[47] br[47] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_50 
+ bl[48] br[48] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_51 
+ bl[49] br[49] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_52 
+ bl[50] br[50] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_53 
+ bl[51] br[51] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_54 
+ bl[52] br[52] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_55 
+ bl[53] br[53] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_56 
+ bl[54] br[54] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_57 
+ bl[55] br[55] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_58 
+ bl[56] br[56] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_59 
+ bl[57] br[57] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_60 
+ bl[58] br[58] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_61 
+ bl[59] br[59] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_62 
+ bl[60] br[60] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_63 
+ bl[61] br[61] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_64 
+ bl[62] br[62] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_65 
+ bl[63] br[63] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_66 
+ bl[64] br[64] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_67 
+ bl[65] br[65] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_68 
+ bl[66] br[66] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_69 
+ bl[67] br[67] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_70 
+ bl[68] br[68] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_71 
+ bl[69] br[69] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_72 
+ bl[70] br[70] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_73 
+ bl[71] br[71] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_74 
+ bl[72] br[72] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_75 
+ bl[73] br[73] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_76 
+ bl[74] br[74] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_77 
+ bl[75] br[75] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_78 
+ bl[76] br[76] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_79 
+ bl[77] br[77] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_80 
+ bl[78] br[78] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_81 
+ bl[79] br[79] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_82 
+ bl[80] br[80] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_83 
+ bl[81] br[81] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_84 
+ bl[82] br[82] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_85 
+ bl[83] br[83] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_86 
+ bl[84] br[84] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_87 
+ bl[85] br[85] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_88 
+ bl[86] br[86] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_89 
+ bl[87] br[87] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_90 
+ bl[88] br[88] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_91 
+ bl[89] br[89] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_92 
+ bl[90] br[90] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_93 
+ bl[91] br[91] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_94 
+ bl[92] br[92] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_95 
+ bl[93] br[93] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_96 
+ bl[94] br[94] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_97 
+ bl[95] br[95] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_98 
+ bl[96] br[96] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_99 
+ bl[97] br[97] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_100 
+ bl[98] br[98] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_101 
+ bl[99] br[99] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_102 
+ bl[100] br[100] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_103 
+ bl[101] br[101] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_104 
+ bl[102] br[102] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_105 
+ bl[103] br[103] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_106 
+ bl[104] br[104] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_107 
+ bl[105] br[105] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_108 
+ bl[106] br[106] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_109 
+ bl[107] br[107] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_110 
+ bl[108] br[108] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_111 
+ bl[109] br[109] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_112 
+ bl[110] br[110] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_113 
+ bl[111] br[111] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_114 
+ bl[112] br[112] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_115 
+ bl[113] br[113] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_116 
+ bl[114] br[114] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_117 
+ bl[115] br[115] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_118 
+ bl[116] br[116] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_119 
+ bl[117] br[117] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_120 
+ bl[118] br[118] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_121 
+ bl[119] br[119] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_122 
+ bl[120] br[120] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_123 
+ bl[121] br[121] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_124 
+ bl[122] br[122] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_125 
+ bl[123] br[123] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_126 
+ bl[124] br[124] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_127 
+ bl[125] br[125] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_128 
+ bl[126] br[126] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_129 
+ bl[127] br[127] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_130 
+ vdd vdd vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_131 
+ vdd vdd vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_0 
+ vdd vdd vss vdd vpb vnb wl[47] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_49_1 
+ rbl rbr vss vdd vpb vnb wl[47] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_49_2 
+ bl[0] br[0] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_3 
+ bl[1] br[1] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_4 
+ bl[2] br[2] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_5 
+ bl[3] br[3] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_6 
+ bl[4] br[4] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_7 
+ bl[5] br[5] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_8 
+ bl[6] br[6] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_9 
+ bl[7] br[7] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_10 
+ bl[8] br[8] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_11 
+ bl[9] br[9] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_12 
+ bl[10] br[10] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_13 
+ bl[11] br[11] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_14 
+ bl[12] br[12] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_15 
+ bl[13] br[13] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_16 
+ bl[14] br[14] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_17 
+ bl[15] br[15] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_18 
+ bl[16] br[16] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_19 
+ bl[17] br[17] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_20 
+ bl[18] br[18] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_21 
+ bl[19] br[19] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_22 
+ bl[20] br[20] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_23 
+ bl[21] br[21] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_24 
+ bl[22] br[22] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_25 
+ bl[23] br[23] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_26 
+ bl[24] br[24] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_27 
+ bl[25] br[25] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_28 
+ bl[26] br[26] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_29 
+ bl[27] br[27] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_30 
+ bl[28] br[28] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_31 
+ bl[29] br[29] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_32 
+ bl[30] br[30] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_33 
+ bl[31] br[31] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_34 
+ bl[32] br[32] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_35 
+ bl[33] br[33] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_36 
+ bl[34] br[34] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_37 
+ bl[35] br[35] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_38 
+ bl[36] br[36] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_39 
+ bl[37] br[37] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_40 
+ bl[38] br[38] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_41 
+ bl[39] br[39] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_42 
+ bl[40] br[40] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_43 
+ bl[41] br[41] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_44 
+ bl[42] br[42] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_45 
+ bl[43] br[43] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_46 
+ bl[44] br[44] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_47 
+ bl[45] br[45] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_48 
+ bl[46] br[46] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_49 
+ bl[47] br[47] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_50 
+ bl[48] br[48] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_51 
+ bl[49] br[49] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_52 
+ bl[50] br[50] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_53 
+ bl[51] br[51] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_54 
+ bl[52] br[52] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_55 
+ bl[53] br[53] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_56 
+ bl[54] br[54] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_57 
+ bl[55] br[55] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_58 
+ bl[56] br[56] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_59 
+ bl[57] br[57] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_60 
+ bl[58] br[58] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_61 
+ bl[59] br[59] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_62 
+ bl[60] br[60] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_63 
+ bl[61] br[61] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_64 
+ bl[62] br[62] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_65 
+ bl[63] br[63] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_66 
+ bl[64] br[64] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_67 
+ bl[65] br[65] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_68 
+ bl[66] br[66] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_69 
+ bl[67] br[67] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_70 
+ bl[68] br[68] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_71 
+ bl[69] br[69] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_72 
+ bl[70] br[70] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_73 
+ bl[71] br[71] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_74 
+ bl[72] br[72] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_75 
+ bl[73] br[73] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_76 
+ bl[74] br[74] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_77 
+ bl[75] br[75] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_78 
+ bl[76] br[76] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_79 
+ bl[77] br[77] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_80 
+ bl[78] br[78] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_81 
+ bl[79] br[79] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_82 
+ bl[80] br[80] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_83 
+ bl[81] br[81] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_84 
+ bl[82] br[82] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_85 
+ bl[83] br[83] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_86 
+ bl[84] br[84] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_87 
+ bl[85] br[85] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_88 
+ bl[86] br[86] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_89 
+ bl[87] br[87] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_90 
+ bl[88] br[88] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_91 
+ bl[89] br[89] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_92 
+ bl[90] br[90] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_93 
+ bl[91] br[91] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_94 
+ bl[92] br[92] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_95 
+ bl[93] br[93] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_96 
+ bl[94] br[94] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_97 
+ bl[95] br[95] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_98 
+ bl[96] br[96] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_99 
+ bl[97] br[97] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_100 
+ bl[98] br[98] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_101 
+ bl[99] br[99] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_102 
+ bl[100] br[100] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_103 
+ bl[101] br[101] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_104 
+ bl[102] br[102] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_105 
+ bl[103] br[103] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_106 
+ bl[104] br[104] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_107 
+ bl[105] br[105] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_108 
+ bl[106] br[106] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_109 
+ bl[107] br[107] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_110 
+ bl[108] br[108] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_111 
+ bl[109] br[109] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_112 
+ bl[110] br[110] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_113 
+ bl[111] br[111] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_114 
+ bl[112] br[112] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_115 
+ bl[113] br[113] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_116 
+ bl[114] br[114] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_117 
+ bl[115] br[115] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_118 
+ bl[116] br[116] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_119 
+ bl[117] br[117] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_120 
+ bl[118] br[118] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_121 
+ bl[119] br[119] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_122 
+ bl[120] br[120] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_123 
+ bl[121] br[121] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_124 
+ bl[122] br[122] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_125 
+ bl[123] br[123] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_126 
+ bl[124] br[124] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_127 
+ bl[125] br[125] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_128 
+ bl[126] br[126] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_129 
+ bl[127] br[127] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_130 
+ vdd vdd vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_131 
+ vdd vdd vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_0 
+ vdd vdd vss vdd vpb vnb wl[48] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_50_1 
+ rbl rbr vss vdd vpb vnb wl[48] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_50_2 
+ bl[0] br[0] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_3 
+ bl[1] br[1] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_4 
+ bl[2] br[2] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_5 
+ bl[3] br[3] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_6 
+ bl[4] br[4] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_7 
+ bl[5] br[5] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_8 
+ bl[6] br[6] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_9 
+ bl[7] br[7] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_10 
+ bl[8] br[8] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_11 
+ bl[9] br[9] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_12 
+ bl[10] br[10] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_13 
+ bl[11] br[11] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_14 
+ bl[12] br[12] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_15 
+ bl[13] br[13] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_16 
+ bl[14] br[14] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_17 
+ bl[15] br[15] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_18 
+ bl[16] br[16] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_19 
+ bl[17] br[17] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_20 
+ bl[18] br[18] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_21 
+ bl[19] br[19] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_22 
+ bl[20] br[20] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_23 
+ bl[21] br[21] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_24 
+ bl[22] br[22] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_25 
+ bl[23] br[23] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_26 
+ bl[24] br[24] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_27 
+ bl[25] br[25] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_28 
+ bl[26] br[26] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_29 
+ bl[27] br[27] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_30 
+ bl[28] br[28] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_31 
+ bl[29] br[29] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_32 
+ bl[30] br[30] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_33 
+ bl[31] br[31] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_34 
+ bl[32] br[32] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_35 
+ bl[33] br[33] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_36 
+ bl[34] br[34] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_37 
+ bl[35] br[35] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_38 
+ bl[36] br[36] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_39 
+ bl[37] br[37] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_40 
+ bl[38] br[38] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_41 
+ bl[39] br[39] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_42 
+ bl[40] br[40] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_43 
+ bl[41] br[41] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_44 
+ bl[42] br[42] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_45 
+ bl[43] br[43] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_46 
+ bl[44] br[44] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_47 
+ bl[45] br[45] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_48 
+ bl[46] br[46] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_49 
+ bl[47] br[47] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_50 
+ bl[48] br[48] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_51 
+ bl[49] br[49] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_52 
+ bl[50] br[50] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_53 
+ bl[51] br[51] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_54 
+ bl[52] br[52] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_55 
+ bl[53] br[53] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_56 
+ bl[54] br[54] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_57 
+ bl[55] br[55] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_58 
+ bl[56] br[56] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_59 
+ bl[57] br[57] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_60 
+ bl[58] br[58] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_61 
+ bl[59] br[59] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_62 
+ bl[60] br[60] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_63 
+ bl[61] br[61] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_64 
+ bl[62] br[62] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_65 
+ bl[63] br[63] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_66 
+ bl[64] br[64] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_67 
+ bl[65] br[65] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_68 
+ bl[66] br[66] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_69 
+ bl[67] br[67] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_70 
+ bl[68] br[68] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_71 
+ bl[69] br[69] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_72 
+ bl[70] br[70] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_73 
+ bl[71] br[71] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_74 
+ bl[72] br[72] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_75 
+ bl[73] br[73] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_76 
+ bl[74] br[74] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_77 
+ bl[75] br[75] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_78 
+ bl[76] br[76] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_79 
+ bl[77] br[77] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_80 
+ bl[78] br[78] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_81 
+ bl[79] br[79] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_82 
+ bl[80] br[80] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_83 
+ bl[81] br[81] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_84 
+ bl[82] br[82] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_85 
+ bl[83] br[83] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_86 
+ bl[84] br[84] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_87 
+ bl[85] br[85] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_88 
+ bl[86] br[86] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_89 
+ bl[87] br[87] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_90 
+ bl[88] br[88] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_91 
+ bl[89] br[89] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_92 
+ bl[90] br[90] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_93 
+ bl[91] br[91] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_94 
+ bl[92] br[92] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_95 
+ bl[93] br[93] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_96 
+ bl[94] br[94] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_97 
+ bl[95] br[95] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_98 
+ bl[96] br[96] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_99 
+ bl[97] br[97] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_100 
+ bl[98] br[98] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_101 
+ bl[99] br[99] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_102 
+ bl[100] br[100] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_103 
+ bl[101] br[101] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_104 
+ bl[102] br[102] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_105 
+ bl[103] br[103] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_106 
+ bl[104] br[104] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_107 
+ bl[105] br[105] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_108 
+ bl[106] br[106] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_109 
+ bl[107] br[107] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_110 
+ bl[108] br[108] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_111 
+ bl[109] br[109] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_112 
+ bl[110] br[110] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_113 
+ bl[111] br[111] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_114 
+ bl[112] br[112] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_115 
+ bl[113] br[113] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_116 
+ bl[114] br[114] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_117 
+ bl[115] br[115] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_118 
+ bl[116] br[116] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_119 
+ bl[117] br[117] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_120 
+ bl[118] br[118] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_121 
+ bl[119] br[119] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_122 
+ bl[120] br[120] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_123 
+ bl[121] br[121] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_124 
+ bl[122] br[122] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_125 
+ bl[123] br[123] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_126 
+ bl[124] br[124] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_127 
+ bl[125] br[125] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_128 
+ bl[126] br[126] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_129 
+ bl[127] br[127] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_130 
+ vdd vdd vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_131 
+ vdd vdd vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_0 
+ vdd vdd vss vdd vpb vnb wl[49] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_51_1 
+ rbl rbr vss vdd vpb vnb wl[49] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_51_2 
+ bl[0] br[0] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_3 
+ bl[1] br[1] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_4 
+ bl[2] br[2] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_5 
+ bl[3] br[3] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_6 
+ bl[4] br[4] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_7 
+ bl[5] br[5] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_8 
+ bl[6] br[6] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_9 
+ bl[7] br[7] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_10 
+ bl[8] br[8] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_11 
+ bl[9] br[9] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_12 
+ bl[10] br[10] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_13 
+ bl[11] br[11] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_14 
+ bl[12] br[12] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_15 
+ bl[13] br[13] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_16 
+ bl[14] br[14] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_17 
+ bl[15] br[15] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_18 
+ bl[16] br[16] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_19 
+ bl[17] br[17] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_20 
+ bl[18] br[18] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_21 
+ bl[19] br[19] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_22 
+ bl[20] br[20] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_23 
+ bl[21] br[21] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_24 
+ bl[22] br[22] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_25 
+ bl[23] br[23] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_26 
+ bl[24] br[24] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_27 
+ bl[25] br[25] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_28 
+ bl[26] br[26] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_29 
+ bl[27] br[27] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_30 
+ bl[28] br[28] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_31 
+ bl[29] br[29] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_32 
+ bl[30] br[30] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_33 
+ bl[31] br[31] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_34 
+ bl[32] br[32] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_35 
+ bl[33] br[33] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_36 
+ bl[34] br[34] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_37 
+ bl[35] br[35] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_38 
+ bl[36] br[36] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_39 
+ bl[37] br[37] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_40 
+ bl[38] br[38] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_41 
+ bl[39] br[39] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_42 
+ bl[40] br[40] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_43 
+ bl[41] br[41] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_44 
+ bl[42] br[42] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_45 
+ bl[43] br[43] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_46 
+ bl[44] br[44] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_47 
+ bl[45] br[45] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_48 
+ bl[46] br[46] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_49 
+ bl[47] br[47] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_50 
+ bl[48] br[48] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_51 
+ bl[49] br[49] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_52 
+ bl[50] br[50] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_53 
+ bl[51] br[51] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_54 
+ bl[52] br[52] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_55 
+ bl[53] br[53] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_56 
+ bl[54] br[54] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_57 
+ bl[55] br[55] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_58 
+ bl[56] br[56] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_59 
+ bl[57] br[57] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_60 
+ bl[58] br[58] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_61 
+ bl[59] br[59] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_62 
+ bl[60] br[60] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_63 
+ bl[61] br[61] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_64 
+ bl[62] br[62] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_65 
+ bl[63] br[63] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_66 
+ bl[64] br[64] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_67 
+ bl[65] br[65] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_68 
+ bl[66] br[66] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_69 
+ bl[67] br[67] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_70 
+ bl[68] br[68] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_71 
+ bl[69] br[69] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_72 
+ bl[70] br[70] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_73 
+ bl[71] br[71] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_74 
+ bl[72] br[72] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_75 
+ bl[73] br[73] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_76 
+ bl[74] br[74] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_77 
+ bl[75] br[75] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_78 
+ bl[76] br[76] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_79 
+ bl[77] br[77] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_80 
+ bl[78] br[78] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_81 
+ bl[79] br[79] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_82 
+ bl[80] br[80] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_83 
+ bl[81] br[81] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_84 
+ bl[82] br[82] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_85 
+ bl[83] br[83] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_86 
+ bl[84] br[84] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_87 
+ bl[85] br[85] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_88 
+ bl[86] br[86] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_89 
+ bl[87] br[87] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_90 
+ bl[88] br[88] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_91 
+ bl[89] br[89] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_92 
+ bl[90] br[90] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_93 
+ bl[91] br[91] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_94 
+ bl[92] br[92] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_95 
+ bl[93] br[93] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_96 
+ bl[94] br[94] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_97 
+ bl[95] br[95] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_98 
+ bl[96] br[96] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_99 
+ bl[97] br[97] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_100 
+ bl[98] br[98] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_101 
+ bl[99] br[99] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_102 
+ bl[100] br[100] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_103 
+ bl[101] br[101] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_104 
+ bl[102] br[102] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_105 
+ bl[103] br[103] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_106 
+ bl[104] br[104] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_107 
+ bl[105] br[105] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_108 
+ bl[106] br[106] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_109 
+ bl[107] br[107] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_110 
+ bl[108] br[108] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_111 
+ bl[109] br[109] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_112 
+ bl[110] br[110] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_113 
+ bl[111] br[111] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_114 
+ bl[112] br[112] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_115 
+ bl[113] br[113] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_116 
+ bl[114] br[114] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_117 
+ bl[115] br[115] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_118 
+ bl[116] br[116] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_119 
+ bl[117] br[117] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_120 
+ bl[118] br[118] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_121 
+ bl[119] br[119] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_122 
+ bl[120] br[120] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_123 
+ bl[121] br[121] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_124 
+ bl[122] br[122] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_125 
+ bl[123] br[123] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_126 
+ bl[124] br[124] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_127 
+ bl[125] br[125] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_128 
+ bl[126] br[126] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_129 
+ bl[127] br[127] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_130 
+ vdd vdd vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_131 
+ vdd vdd vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_0 
+ vdd vdd vss vdd vpb vnb wl[50] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_52_1 
+ rbl rbr vss vdd vpb vnb wl[50] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_52_2 
+ bl[0] br[0] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_3 
+ bl[1] br[1] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_4 
+ bl[2] br[2] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_5 
+ bl[3] br[3] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_6 
+ bl[4] br[4] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_7 
+ bl[5] br[5] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_8 
+ bl[6] br[6] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_9 
+ bl[7] br[7] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_10 
+ bl[8] br[8] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_11 
+ bl[9] br[9] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_12 
+ bl[10] br[10] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_13 
+ bl[11] br[11] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_14 
+ bl[12] br[12] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_15 
+ bl[13] br[13] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_16 
+ bl[14] br[14] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_17 
+ bl[15] br[15] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_18 
+ bl[16] br[16] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_19 
+ bl[17] br[17] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_20 
+ bl[18] br[18] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_21 
+ bl[19] br[19] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_22 
+ bl[20] br[20] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_23 
+ bl[21] br[21] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_24 
+ bl[22] br[22] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_25 
+ bl[23] br[23] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_26 
+ bl[24] br[24] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_27 
+ bl[25] br[25] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_28 
+ bl[26] br[26] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_29 
+ bl[27] br[27] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_30 
+ bl[28] br[28] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_31 
+ bl[29] br[29] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_32 
+ bl[30] br[30] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_33 
+ bl[31] br[31] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_34 
+ bl[32] br[32] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_35 
+ bl[33] br[33] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_36 
+ bl[34] br[34] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_37 
+ bl[35] br[35] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_38 
+ bl[36] br[36] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_39 
+ bl[37] br[37] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_40 
+ bl[38] br[38] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_41 
+ bl[39] br[39] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_42 
+ bl[40] br[40] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_43 
+ bl[41] br[41] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_44 
+ bl[42] br[42] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_45 
+ bl[43] br[43] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_46 
+ bl[44] br[44] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_47 
+ bl[45] br[45] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_48 
+ bl[46] br[46] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_49 
+ bl[47] br[47] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_50 
+ bl[48] br[48] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_51 
+ bl[49] br[49] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_52 
+ bl[50] br[50] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_53 
+ bl[51] br[51] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_54 
+ bl[52] br[52] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_55 
+ bl[53] br[53] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_56 
+ bl[54] br[54] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_57 
+ bl[55] br[55] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_58 
+ bl[56] br[56] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_59 
+ bl[57] br[57] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_60 
+ bl[58] br[58] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_61 
+ bl[59] br[59] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_62 
+ bl[60] br[60] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_63 
+ bl[61] br[61] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_64 
+ bl[62] br[62] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_65 
+ bl[63] br[63] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_66 
+ bl[64] br[64] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_67 
+ bl[65] br[65] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_68 
+ bl[66] br[66] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_69 
+ bl[67] br[67] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_70 
+ bl[68] br[68] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_71 
+ bl[69] br[69] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_72 
+ bl[70] br[70] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_73 
+ bl[71] br[71] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_74 
+ bl[72] br[72] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_75 
+ bl[73] br[73] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_76 
+ bl[74] br[74] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_77 
+ bl[75] br[75] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_78 
+ bl[76] br[76] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_79 
+ bl[77] br[77] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_80 
+ bl[78] br[78] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_81 
+ bl[79] br[79] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_82 
+ bl[80] br[80] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_83 
+ bl[81] br[81] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_84 
+ bl[82] br[82] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_85 
+ bl[83] br[83] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_86 
+ bl[84] br[84] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_87 
+ bl[85] br[85] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_88 
+ bl[86] br[86] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_89 
+ bl[87] br[87] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_90 
+ bl[88] br[88] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_91 
+ bl[89] br[89] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_92 
+ bl[90] br[90] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_93 
+ bl[91] br[91] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_94 
+ bl[92] br[92] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_95 
+ bl[93] br[93] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_96 
+ bl[94] br[94] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_97 
+ bl[95] br[95] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_98 
+ bl[96] br[96] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_99 
+ bl[97] br[97] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_100 
+ bl[98] br[98] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_101 
+ bl[99] br[99] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_102 
+ bl[100] br[100] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_103 
+ bl[101] br[101] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_104 
+ bl[102] br[102] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_105 
+ bl[103] br[103] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_106 
+ bl[104] br[104] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_107 
+ bl[105] br[105] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_108 
+ bl[106] br[106] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_109 
+ bl[107] br[107] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_110 
+ bl[108] br[108] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_111 
+ bl[109] br[109] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_112 
+ bl[110] br[110] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_113 
+ bl[111] br[111] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_114 
+ bl[112] br[112] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_115 
+ bl[113] br[113] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_116 
+ bl[114] br[114] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_117 
+ bl[115] br[115] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_118 
+ bl[116] br[116] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_119 
+ bl[117] br[117] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_120 
+ bl[118] br[118] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_121 
+ bl[119] br[119] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_122 
+ bl[120] br[120] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_123 
+ bl[121] br[121] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_124 
+ bl[122] br[122] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_125 
+ bl[123] br[123] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_126 
+ bl[124] br[124] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_127 
+ bl[125] br[125] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_128 
+ bl[126] br[126] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_129 
+ bl[127] br[127] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_130 
+ vdd vdd vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_131 
+ vdd vdd vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_0 
+ vdd vdd vss vdd vpb vnb wl[51] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_53_1 
+ rbl rbr vss vdd vpb vnb wl[51] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_53_2 
+ bl[0] br[0] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_3 
+ bl[1] br[1] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_4 
+ bl[2] br[2] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_5 
+ bl[3] br[3] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_6 
+ bl[4] br[4] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_7 
+ bl[5] br[5] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_8 
+ bl[6] br[6] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_9 
+ bl[7] br[7] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_10 
+ bl[8] br[8] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_11 
+ bl[9] br[9] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_12 
+ bl[10] br[10] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_13 
+ bl[11] br[11] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_14 
+ bl[12] br[12] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_15 
+ bl[13] br[13] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_16 
+ bl[14] br[14] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_17 
+ bl[15] br[15] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_18 
+ bl[16] br[16] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_19 
+ bl[17] br[17] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_20 
+ bl[18] br[18] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_21 
+ bl[19] br[19] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_22 
+ bl[20] br[20] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_23 
+ bl[21] br[21] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_24 
+ bl[22] br[22] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_25 
+ bl[23] br[23] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_26 
+ bl[24] br[24] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_27 
+ bl[25] br[25] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_28 
+ bl[26] br[26] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_29 
+ bl[27] br[27] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_30 
+ bl[28] br[28] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_31 
+ bl[29] br[29] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_32 
+ bl[30] br[30] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_33 
+ bl[31] br[31] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_34 
+ bl[32] br[32] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_35 
+ bl[33] br[33] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_36 
+ bl[34] br[34] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_37 
+ bl[35] br[35] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_38 
+ bl[36] br[36] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_39 
+ bl[37] br[37] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_40 
+ bl[38] br[38] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_41 
+ bl[39] br[39] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_42 
+ bl[40] br[40] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_43 
+ bl[41] br[41] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_44 
+ bl[42] br[42] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_45 
+ bl[43] br[43] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_46 
+ bl[44] br[44] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_47 
+ bl[45] br[45] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_48 
+ bl[46] br[46] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_49 
+ bl[47] br[47] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_50 
+ bl[48] br[48] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_51 
+ bl[49] br[49] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_52 
+ bl[50] br[50] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_53 
+ bl[51] br[51] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_54 
+ bl[52] br[52] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_55 
+ bl[53] br[53] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_56 
+ bl[54] br[54] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_57 
+ bl[55] br[55] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_58 
+ bl[56] br[56] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_59 
+ bl[57] br[57] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_60 
+ bl[58] br[58] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_61 
+ bl[59] br[59] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_62 
+ bl[60] br[60] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_63 
+ bl[61] br[61] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_64 
+ bl[62] br[62] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_65 
+ bl[63] br[63] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_66 
+ bl[64] br[64] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_67 
+ bl[65] br[65] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_68 
+ bl[66] br[66] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_69 
+ bl[67] br[67] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_70 
+ bl[68] br[68] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_71 
+ bl[69] br[69] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_72 
+ bl[70] br[70] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_73 
+ bl[71] br[71] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_74 
+ bl[72] br[72] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_75 
+ bl[73] br[73] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_76 
+ bl[74] br[74] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_77 
+ bl[75] br[75] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_78 
+ bl[76] br[76] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_79 
+ bl[77] br[77] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_80 
+ bl[78] br[78] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_81 
+ bl[79] br[79] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_82 
+ bl[80] br[80] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_83 
+ bl[81] br[81] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_84 
+ bl[82] br[82] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_85 
+ bl[83] br[83] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_86 
+ bl[84] br[84] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_87 
+ bl[85] br[85] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_88 
+ bl[86] br[86] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_89 
+ bl[87] br[87] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_90 
+ bl[88] br[88] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_91 
+ bl[89] br[89] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_92 
+ bl[90] br[90] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_93 
+ bl[91] br[91] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_94 
+ bl[92] br[92] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_95 
+ bl[93] br[93] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_96 
+ bl[94] br[94] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_97 
+ bl[95] br[95] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_98 
+ bl[96] br[96] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_99 
+ bl[97] br[97] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_100 
+ bl[98] br[98] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_101 
+ bl[99] br[99] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_102 
+ bl[100] br[100] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_103 
+ bl[101] br[101] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_104 
+ bl[102] br[102] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_105 
+ bl[103] br[103] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_106 
+ bl[104] br[104] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_107 
+ bl[105] br[105] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_108 
+ bl[106] br[106] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_109 
+ bl[107] br[107] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_110 
+ bl[108] br[108] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_111 
+ bl[109] br[109] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_112 
+ bl[110] br[110] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_113 
+ bl[111] br[111] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_114 
+ bl[112] br[112] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_115 
+ bl[113] br[113] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_116 
+ bl[114] br[114] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_117 
+ bl[115] br[115] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_118 
+ bl[116] br[116] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_119 
+ bl[117] br[117] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_120 
+ bl[118] br[118] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_121 
+ bl[119] br[119] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_122 
+ bl[120] br[120] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_123 
+ bl[121] br[121] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_124 
+ bl[122] br[122] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_125 
+ bl[123] br[123] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_126 
+ bl[124] br[124] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_127 
+ bl[125] br[125] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_128 
+ bl[126] br[126] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_129 
+ bl[127] br[127] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_130 
+ vdd vdd vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_131 
+ vdd vdd vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_0 
+ vdd vdd vss vdd vpb vnb wl[52] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_54_1 
+ rbl rbr vss vdd vpb vnb wl[52] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_54_2 
+ bl[0] br[0] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_3 
+ bl[1] br[1] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_4 
+ bl[2] br[2] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_5 
+ bl[3] br[3] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_6 
+ bl[4] br[4] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_7 
+ bl[5] br[5] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_8 
+ bl[6] br[6] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_9 
+ bl[7] br[7] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_10 
+ bl[8] br[8] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_11 
+ bl[9] br[9] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_12 
+ bl[10] br[10] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_13 
+ bl[11] br[11] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_14 
+ bl[12] br[12] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_15 
+ bl[13] br[13] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_16 
+ bl[14] br[14] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_17 
+ bl[15] br[15] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_18 
+ bl[16] br[16] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_19 
+ bl[17] br[17] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_20 
+ bl[18] br[18] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_21 
+ bl[19] br[19] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_22 
+ bl[20] br[20] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_23 
+ bl[21] br[21] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_24 
+ bl[22] br[22] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_25 
+ bl[23] br[23] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_26 
+ bl[24] br[24] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_27 
+ bl[25] br[25] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_28 
+ bl[26] br[26] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_29 
+ bl[27] br[27] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_30 
+ bl[28] br[28] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_31 
+ bl[29] br[29] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_32 
+ bl[30] br[30] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_33 
+ bl[31] br[31] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_34 
+ bl[32] br[32] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_35 
+ bl[33] br[33] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_36 
+ bl[34] br[34] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_37 
+ bl[35] br[35] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_38 
+ bl[36] br[36] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_39 
+ bl[37] br[37] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_40 
+ bl[38] br[38] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_41 
+ bl[39] br[39] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_42 
+ bl[40] br[40] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_43 
+ bl[41] br[41] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_44 
+ bl[42] br[42] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_45 
+ bl[43] br[43] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_46 
+ bl[44] br[44] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_47 
+ bl[45] br[45] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_48 
+ bl[46] br[46] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_49 
+ bl[47] br[47] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_50 
+ bl[48] br[48] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_51 
+ bl[49] br[49] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_52 
+ bl[50] br[50] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_53 
+ bl[51] br[51] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_54 
+ bl[52] br[52] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_55 
+ bl[53] br[53] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_56 
+ bl[54] br[54] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_57 
+ bl[55] br[55] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_58 
+ bl[56] br[56] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_59 
+ bl[57] br[57] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_60 
+ bl[58] br[58] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_61 
+ bl[59] br[59] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_62 
+ bl[60] br[60] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_63 
+ bl[61] br[61] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_64 
+ bl[62] br[62] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_65 
+ bl[63] br[63] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_66 
+ bl[64] br[64] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_67 
+ bl[65] br[65] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_68 
+ bl[66] br[66] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_69 
+ bl[67] br[67] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_70 
+ bl[68] br[68] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_71 
+ bl[69] br[69] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_72 
+ bl[70] br[70] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_73 
+ bl[71] br[71] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_74 
+ bl[72] br[72] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_75 
+ bl[73] br[73] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_76 
+ bl[74] br[74] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_77 
+ bl[75] br[75] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_78 
+ bl[76] br[76] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_79 
+ bl[77] br[77] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_80 
+ bl[78] br[78] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_81 
+ bl[79] br[79] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_82 
+ bl[80] br[80] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_83 
+ bl[81] br[81] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_84 
+ bl[82] br[82] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_85 
+ bl[83] br[83] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_86 
+ bl[84] br[84] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_87 
+ bl[85] br[85] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_88 
+ bl[86] br[86] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_89 
+ bl[87] br[87] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_90 
+ bl[88] br[88] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_91 
+ bl[89] br[89] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_92 
+ bl[90] br[90] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_93 
+ bl[91] br[91] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_94 
+ bl[92] br[92] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_95 
+ bl[93] br[93] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_96 
+ bl[94] br[94] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_97 
+ bl[95] br[95] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_98 
+ bl[96] br[96] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_99 
+ bl[97] br[97] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_100 
+ bl[98] br[98] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_101 
+ bl[99] br[99] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_102 
+ bl[100] br[100] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_103 
+ bl[101] br[101] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_104 
+ bl[102] br[102] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_105 
+ bl[103] br[103] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_106 
+ bl[104] br[104] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_107 
+ bl[105] br[105] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_108 
+ bl[106] br[106] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_109 
+ bl[107] br[107] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_110 
+ bl[108] br[108] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_111 
+ bl[109] br[109] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_112 
+ bl[110] br[110] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_113 
+ bl[111] br[111] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_114 
+ bl[112] br[112] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_115 
+ bl[113] br[113] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_116 
+ bl[114] br[114] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_117 
+ bl[115] br[115] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_118 
+ bl[116] br[116] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_119 
+ bl[117] br[117] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_120 
+ bl[118] br[118] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_121 
+ bl[119] br[119] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_122 
+ bl[120] br[120] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_123 
+ bl[121] br[121] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_124 
+ bl[122] br[122] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_125 
+ bl[123] br[123] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_126 
+ bl[124] br[124] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_127 
+ bl[125] br[125] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_128 
+ bl[126] br[126] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_129 
+ bl[127] br[127] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_130 
+ vdd vdd vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_131 
+ vdd vdd vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_0 
+ vdd vdd vss vdd vpb vnb wl[53] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_55_1 
+ rbl rbr vss vdd vpb vnb wl[53] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_55_2 
+ bl[0] br[0] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_3 
+ bl[1] br[1] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_4 
+ bl[2] br[2] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_5 
+ bl[3] br[3] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_6 
+ bl[4] br[4] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_7 
+ bl[5] br[5] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_8 
+ bl[6] br[6] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_9 
+ bl[7] br[7] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_10 
+ bl[8] br[8] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_11 
+ bl[9] br[9] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_12 
+ bl[10] br[10] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_13 
+ bl[11] br[11] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_14 
+ bl[12] br[12] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_15 
+ bl[13] br[13] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_16 
+ bl[14] br[14] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_17 
+ bl[15] br[15] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_18 
+ bl[16] br[16] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_19 
+ bl[17] br[17] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_20 
+ bl[18] br[18] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_21 
+ bl[19] br[19] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_22 
+ bl[20] br[20] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_23 
+ bl[21] br[21] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_24 
+ bl[22] br[22] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_25 
+ bl[23] br[23] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_26 
+ bl[24] br[24] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_27 
+ bl[25] br[25] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_28 
+ bl[26] br[26] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_29 
+ bl[27] br[27] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_30 
+ bl[28] br[28] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_31 
+ bl[29] br[29] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_32 
+ bl[30] br[30] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_33 
+ bl[31] br[31] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_34 
+ bl[32] br[32] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_35 
+ bl[33] br[33] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_36 
+ bl[34] br[34] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_37 
+ bl[35] br[35] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_38 
+ bl[36] br[36] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_39 
+ bl[37] br[37] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_40 
+ bl[38] br[38] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_41 
+ bl[39] br[39] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_42 
+ bl[40] br[40] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_43 
+ bl[41] br[41] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_44 
+ bl[42] br[42] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_45 
+ bl[43] br[43] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_46 
+ bl[44] br[44] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_47 
+ bl[45] br[45] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_48 
+ bl[46] br[46] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_49 
+ bl[47] br[47] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_50 
+ bl[48] br[48] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_51 
+ bl[49] br[49] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_52 
+ bl[50] br[50] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_53 
+ bl[51] br[51] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_54 
+ bl[52] br[52] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_55 
+ bl[53] br[53] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_56 
+ bl[54] br[54] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_57 
+ bl[55] br[55] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_58 
+ bl[56] br[56] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_59 
+ bl[57] br[57] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_60 
+ bl[58] br[58] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_61 
+ bl[59] br[59] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_62 
+ bl[60] br[60] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_63 
+ bl[61] br[61] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_64 
+ bl[62] br[62] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_65 
+ bl[63] br[63] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_66 
+ bl[64] br[64] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_67 
+ bl[65] br[65] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_68 
+ bl[66] br[66] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_69 
+ bl[67] br[67] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_70 
+ bl[68] br[68] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_71 
+ bl[69] br[69] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_72 
+ bl[70] br[70] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_73 
+ bl[71] br[71] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_74 
+ bl[72] br[72] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_75 
+ bl[73] br[73] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_76 
+ bl[74] br[74] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_77 
+ bl[75] br[75] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_78 
+ bl[76] br[76] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_79 
+ bl[77] br[77] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_80 
+ bl[78] br[78] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_81 
+ bl[79] br[79] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_82 
+ bl[80] br[80] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_83 
+ bl[81] br[81] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_84 
+ bl[82] br[82] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_85 
+ bl[83] br[83] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_86 
+ bl[84] br[84] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_87 
+ bl[85] br[85] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_88 
+ bl[86] br[86] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_89 
+ bl[87] br[87] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_90 
+ bl[88] br[88] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_91 
+ bl[89] br[89] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_92 
+ bl[90] br[90] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_93 
+ bl[91] br[91] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_94 
+ bl[92] br[92] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_95 
+ bl[93] br[93] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_96 
+ bl[94] br[94] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_97 
+ bl[95] br[95] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_98 
+ bl[96] br[96] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_99 
+ bl[97] br[97] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_100 
+ bl[98] br[98] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_101 
+ bl[99] br[99] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_102 
+ bl[100] br[100] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_103 
+ bl[101] br[101] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_104 
+ bl[102] br[102] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_105 
+ bl[103] br[103] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_106 
+ bl[104] br[104] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_107 
+ bl[105] br[105] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_108 
+ bl[106] br[106] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_109 
+ bl[107] br[107] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_110 
+ bl[108] br[108] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_111 
+ bl[109] br[109] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_112 
+ bl[110] br[110] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_113 
+ bl[111] br[111] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_114 
+ bl[112] br[112] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_115 
+ bl[113] br[113] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_116 
+ bl[114] br[114] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_117 
+ bl[115] br[115] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_118 
+ bl[116] br[116] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_119 
+ bl[117] br[117] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_120 
+ bl[118] br[118] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_121 
+ bl[119] br[119] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_122 
+ bl[120] br[120] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_123 
+ bl[121] br[121] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_124 
+ bl[122] br[122] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_125 
+ bl[123] br[123] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_126 
+ bl[124] br[124] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_127 
+ bl[125] br[125] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_128 
+ bl[126] br[126] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_129 
+ bl[127] br[127] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_130 
+ vdd vdd vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_131 
+ vdd vdd vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_0 
+ vdd vdd vss vdd vpb vnb wl[54] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_56_1 
+ rbl rbr vss vdd vpb vnb wl[54] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_56_2 
+ bl[0] br[0] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_3 
+ bl[1] br[1] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_4 
+ bl[2] br[2] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_5 
+ bl[3] br[3] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_6 
+ bl[4] br[4] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_7 
+ bl[5] br[5] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_8 
+ bl[6] br[6] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_9 
+ bl[7] br[7] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_10 
+ bl[8] br[8] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_11 
+ bl[9] br[9] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_12 
+ bl[10] br[10] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_13 
+ bl[11] br[11] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_14 
+ bl[12] br[12] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_15 
+ bl[13] br[13] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_16 
+ bl[14] br[14] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_17 
+ bl[15] br[15] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_18 
+ bl[16] br[16] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_19 
+ bl[17] br[17] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_20 
+ bl[18] br[18] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_21 
+ bl[19] br[19] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_22 
+ bl[20] br[20] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_23 
+ bl[21] br[21] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_24 
+ bl[22] br[22] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_25 
+ bl[23] br[23] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_26 
+ bl[24] br[24] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_27 
+ bl[25] br[25] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_28 
+ bl[26] br[26] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_29 
+ bl[27] br[27] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_30 
+ bl[28] br[28] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_31 
+ bl[29] br[29] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_32 
+ bl[30] br[30] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_33 
+ bl[31] br[31] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_34 
+ bl[32] br[32] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_35 
+ bl[33] br[33] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_36 
+ bl[34] br[34] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_37 
+ bl[35] br[35] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_38 
+ bl[36] br[36] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_39 
+ bl[37] br[37] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_40 
+ bl[38] br[38] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_41 
+ bl[39] br[39] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_42 
+ bl[40] br[40] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_43 
+ bl[41] br[41] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_44 
+ bl[42] br[42] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_45 
+ bl[43] br[43] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_46 
+ bl[44] br[44] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_47 
+ bl[45] br[45] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_48 
+ bl[46] br[46] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_49 
+ bl[47] br[47] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_50 
+ bl[48] br[48] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_51 
+ bl[49] br[49] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_52 
+ bl[50] br[50] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_53 
+ bl[51] br[51] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_54 
+ bl[52] br[52] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_55 
+ bl[53] br[53] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_56 
+ bl[54] br[54] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_57 
+ bl[55] br[55] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_58 
+ bl[56] br[56] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_59 
+ bl[57] br[57] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_60 
+ bl[58] br[58] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_61 
+ bl[59] br[59] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_62 
+ bl[60] br[60] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_63 
+ bl[61] br[61] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_64 
+ bl[62] br[62] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_65 
+ bl[63] br[63] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_66 
+ bl[64] br[64] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_67 
+ bl[65] br[65] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_68 
+ bl[66] br[66] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_69 
+ bl[67] br[67] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_70 
+ bl[68] br[68] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_71 
+ bl[69] br[69] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_72 
+ bl[70] br[70] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_73 
+ bl[71] br[71] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_74 
+ bl[72] br[72] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_75 
+ bl[73] br[73] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_76 
+ bl[74] br[74] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_77 
+ bl[75] br[75] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_78 
+ bl[76] br[76] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_79 
+ bl[77] br[77] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_80 
+ bl[78] br[78] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_81 
+ bl[79] br[79] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_82 
+ bl[80] br[80] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_83 
+ bl[81] br[81] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_84 
+ bl[82] br[82] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_85 
+ bl[83] br[83] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_86 
+ bl[84] br[84] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_87 
+ bl[85] br[85] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_88 
+ bl[86] br[86] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_89 
+ bl[87] br[87] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_90 
+ bl[88] br[88] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_91 
+ bl[89] br[89] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_92 
+ bl[90] br[90] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_93 
+ bl[91] br[91] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_94 
+ bl[92] br[92] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_95 
+ bl[93] br[93] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_96 
+ bl[94] br[94] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_97 
+ bl[95] br[95] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_98 
+ bl[96] br[96] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_99 
+ bl[97] br[97] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_100 
+ bl[98] br[98] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_101 
+ bl[99] br[99] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_102 
+ bl[100] br[100] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_103 
+ bl[101] br[101] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_104 
+ bl[102] br[102] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_105 
+ bl[103] br[103] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_106 
+ bl[104] br[104] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_107 
+ bl[105] br[105] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_108 
+ bl[106] br[106] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_109 
+ bl[107] br[107] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_110 
+ bl[108] br[108] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_111 
+ bl[109] br[109] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_112 
+ bl[110] br[110] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_113 
+ bl[111] br[111] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_114 
+ bl[112] br[112] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_115 
+ bl[113] br[113] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_116 
+ bl[114] br[114] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_117 
+ bl[115] br[115] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_118 
+ bl[116] br[116] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_119 
+ bl[117] br[117] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_120 
+ bl[118] br[118] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_121 
+ bl[119] br[119] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_122 
+ bl[120] br[120] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_123 
+ bl[121] br[121] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_124 
+ bl[122] br[122] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_125 
+ bl[123] br[123] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_126 
+ bl[124] br[124] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_127 
+ bl[125] br[125] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_128 
+ bl[126] br[126] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_129 
+ bl[127] br[127] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_130 
+ vdd vdd vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_131 
+ vdd vdd vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_0 
+ vdd vdd vss vdd vpb vnb wl[55] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_57_1 
+ rbl rbr vss vdd vpb vnb wl[55] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_57_2 
+ bl[0] br[0] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_3 
+ bl[1] br[1] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_4 
+ bl[2] br[2] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_5 
+ bl[3] br[3] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_6 
+ bl[4] br[4] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_7 
+ bl[5] br[5] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_8 
+ bl[6] br[6] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_9 
+ bl[7] br[7] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_10 
+ bl[8] br[8] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_11 
+ bl[9] br[9] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_12 
+ bl[10] br[10] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_13 
+ bl[11] br[11] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_14 
+ bl[12] br[12] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_15 
+ bl[13] br[13] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_16 
+ bl[14] br[14] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_17 
+ bl[15] br[15] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_18 
+ bl[16] br[16] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_19 
+ bl[17] br[17] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_20 
+ bl[18] br[18] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_21 
+ bl[19] br[19] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_22 
+ bl[20] br[20] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_23 
+ bl[21] br[21] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_24 
+ bl[22] br[22] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_25 
+ bl[23] br[23] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_26 
+ bl[24] br[24] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_27 
+ bl[25] br[25] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_28 
+ bl[26] br[26] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_29 
+ bl[27] br[27] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_30 
+ bl[28] br[28] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_31 
+ bl[29] br[29] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_32 
+ bl[30] br[30] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_33 
+ bl[31] br[31] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_34 
+ bl[32] br[32] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_35 
+ bl[33] br[33] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_36 
+ bl[34] br[34] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_37 
+ bl[35] br[35] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_38 
+ bl[36] br[36] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_39 
+ bl[37] br[37] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_40 
+ bl[38] br[38] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_41 
+ bl[39] br[39] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_42 
+ bl[40] br[40] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_43 
+ bl[41] br[41] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_44 
+ bl[42] br[42] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_45 
+ bl[43] br[43] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_46 
+ bl[44] br[44] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_47 
+ bl[45] br[45] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_48 
+ bl[46] br[46] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_49 
+ bl[47] br[47] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_50 
+ bl[48] br[48] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_51 
+ bl[49] br[49] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_52 
+ bl[50] br[50] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_53 
+ bl[51] br[51] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_54 
+ bl[52] br[52] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_55 
+ bl[53] br[53] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_56 
+ bl[54] br[54] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_57 
+ bl[55] br[55] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_58 
+ bl[56] br[56] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_59 
+ bl[57] br[57] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_60 
+ bl[58] br[58] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_61 
+ bl[59] br[59] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_62 
+ bl[60] br[60] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_63 
+ bl[61] br[61] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_64 
+ bl[62] br[62] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_65 
+ bl[63] br[63] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_66 
+ bl[64] br[64] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_67 
+ bl[65] br[65] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_68 
+ bl[66] br[66] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_69 
+ bl[67] br[67] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_70 
+ bl[68] br[68] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_71 
+ bl[69] br[69] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_72 
+ bl[70] br[70] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_73 
+ bl[71] br[71] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_74 
+ bl[72] br[72] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_75 
+ bl[73] br[73] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_76 
+ bl[74] br[74] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_77 
+ bl[75] br[75] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_78 
+ bl[76] br[76] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_79 
+ bl[77] br[77] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_80 
+ bl[78] br[78] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_81 
+ bl[79] br[79] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_82 
+ bl[80] br[80] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_83 
+ bl[81] br[81] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_84 
+ bl[82] br[82] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_85 
+ bl[83] br[83] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_86 
+ bl[84] br[84] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_87 
+ bl[85] br[85] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_88 
+ bl[86] br[86] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_89 
+ bl[87] br[87] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_90 
+ bl[88] br[88] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_91 
+ bl[89] br[89] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_92 
+ bl[90] br[90] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_93 
+ bl[91] br[91] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_94 
+ bl[92] br[92] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_95 
+ bl[93] br[93] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_96 
+ bl[94] br[94] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_97 
+ bl[95] br[95] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_98 
+ bl[96] br[96] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_99 
+ bl[97] br[97] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_100 
+ bl[98] br[98] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_101 
+ bl[99] br[99] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_102 
+ bl[100] br[100] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_103 
+ bl[101] br[101] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_104 
+ bl[102] br[102] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_105 
+ bl[103] br[103] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_106 
+ bl[104] br[104] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_107 
+ bl[105] br[105] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_108 
+ bl[106] br[106] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_109 
+ bl[107] br[107] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_110 
+ bl[108] br[108] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_111 
+ bl[109] br[109] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_112 
+ bl[110] br[110] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_113 
+ bl[111] br[111] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_114 
+ bl[112] br[112] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_115 
+ bl[113] br[113] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_116 
+ bl[114] br[114] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_117 
+ bl[115] br[115] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_118 
+ bl[116] br[116] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_119 
+ bl[117] br[117] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_120 
+ bl[118] br[118] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_121 
+ bl[119] br[119] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_122 
+ bl[120] br[120] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_123 
+ bl[121] br[121] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_124 
+ bl[122] br[122] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_125 
+ bl[123] br[123] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_126 
+ bl[124] br[124] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_127 
+ bl[125] br[125] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_128 
+ bl[126] br[126] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_129 
+ bl[127] br[127] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_130 
+ vdd vdd vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_131 
+ vdd vdd vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_0 
+ vdd vdd vss vdd vpb vnb wl[56] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_58_1 
+ rbl rbr vss vdd vpb vnb wl[56] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_58_2 
+ bl[0] br[0] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_3 
+ bl[1] br[1] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_4 
+ bl[2] br[2] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_5 
+ bl[3] br[3] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_6 
+ bl[4] br[4] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_7 
+ bl[5] br[5] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_8 
+ bl[6] br[6] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_9 
+ bl[7] br[7] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_10 
+ bl[8] br[8] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_11 
+ bl[9] br[9] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_12 
+ bl[10] br[10] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_13 
+ bl[11] br[11] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_14 
+ bl[12] br[12] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_15 
+ bl[13] br[13] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_16 
+ bl[14] br[14] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_17 
+ bl[15] br[15] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_18 
+ bl[16] br[16] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_19 
+ bl[17] br[17] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_20 
+ bl[18] br[18] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_21 
+ bl[19] br[19] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_22 
+ bl[20] br[20] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_23 
+ bl[21] br[21] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_24 
+ bl[22] br[22] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_25 
+ bl[23] br[23] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_26 
+ bl[24] br[24] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_27 
+ bl[25] br[25] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_28 
+ bl[26] br[26] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_29 
+ bl[27] br[27] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_30 
+ bl[28] br[28] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_31 
+ bl[29] br[29] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_32 
+ bl[30] br[30] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_33 
+ bl[31] br[31] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_34 
+ bl[32] br[32] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_35 
+ bl[33] br[33] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_36 
+ bl[34] br[34] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_37 
+ bl[35] br[35] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_38 
+ bl[36] br[36] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_39 
+ bl[37] br[37] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_40 
+ bl[38] br[38] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_41 
+ bl[39] br[39] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_42 
+ bl[40] br[40] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_43 
+ bl[41] br[41] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_44 
+ bl[42] br[42] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_45 
+ bl[43] br[43] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_46 
+ bl[44] br[44] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_47 
+ bl[45] br[45] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_48 
+ bl[46] br[46] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_49 
+ bl[47] br[47] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_50 
+ bl[48] br[48] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_51 
+ bl[49] br[49] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_52 
+ bl[50] br[50] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_53 
+ bl[51] br[51] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_54 
+ bl[52] br[52] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_55 
+ bl[53] br[53] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_56 
+ bl[54] br[54] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_57 
+ bl[55] br[55] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_58 
+ bl[56] br[56] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_59 
+ bl[57] br[57] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_60 
+ bl[58] br[58] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_61 
+ bl[59] br[59] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_62 
+ bl[60] br[60] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_63 
+ bl[61] br[61] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_64 
+ bl[62] br[62] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_65 
+ bl[63] br[63] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_66 
+ bl[64] br[64] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_67 
+ bl[65] br[65] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_68 
+ bl[66] br[66] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_69 
+ bl[67] br[67] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_70 
+ bl[68] br[68] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_71 
+ bl[69] br[69] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_72 
+ bl[70] br[70] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_73 
+ bl[71] br[71] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_74 
+ bl[72] br[72] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_75 
+ bl[73] br[73] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_76 
+ bl[74] br[74] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_77 
+ bl[75] br[75] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_78 
+ bl[76] br[76] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_79 
+ bl[77] br[77] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_80 
+ bl[78] br[78] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_81 
+ bl[79] br[79] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_82 
+ bl[80] br[80] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_83 
+ bl[81] br[81] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_84 
+ bl[82] br[82] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_85 
+ bl[83] br[83] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_86 
+ bl[84] br[84] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_87 
+ bl[85] br[85] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_88 
+ bl[86] br[86] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_89 
+ bl[87] br[87] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_90 
+ bl[88] br[88] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_91 
+ bl[89] br[89] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_92 
+ bl[90] br[90] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_93 
+ bl[91] br[91] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_94 
+ bl[92] br[92] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_95 
+ bl[93] br[93] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_96 
+ bl[94] br[94] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_97 
+ bl[95] br[95] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_98 
+ bl[96] br[96] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_99 
+ bl[97] br[97] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_100 
+ bl[98] br[98] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_101 
+ bl[99] br[99] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_102 
+ bl[100] br[100] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_103 
+ bl[101] br[101] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_104 
+ bl[102] br[102] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_105 
+ bl[103] br[103] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_106 
+ bl[104] br[104] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_107 
+ bl[105] br[105] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_108 
+ bl[106] br[106] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_109 
+ bl[107] br[107] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_110 
+ bl[108] br[108] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_111 
+ bl[109] br[109] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_112 
+ bl[110] br[110] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_113 
+ bl[111] br[111] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_114 
+ bl[112] br[112] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_115 
+ bl[113] br[113] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_116 
+ bl[114] br[114] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_117 
+ bl[115] br[115] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_118 
+ bl[116] br[116] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_119 
+ bl[117] br[117] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_120 
+ bl[118] br[118] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_121 
+ bl[119] br[119] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_122 
+ bl[120] br[120] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_123 
+ bl[121] br[121] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_124 
+ bl[122] br[122] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_125 
+ bl[123] br[123] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_126 
+ bl[124] br[124] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_127 
+ bl[125] br[125] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_128 
+ bl[126] br[126] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_129 
+ bl[127] br[127] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_130 
+ vdd vdd vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_131 
+ vdd vdd vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_0 
+ vdd vdd vss vdd vpb vnb wl[57] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_59_1 
+ rbl rbr vss vdd vpb vnb wl[57] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_59_2 
+ bl[0] br[0] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_3 
+ bl[1] br[1] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_4 
+ bl[2] br[2] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_5 
+ bl[3] br[3] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_6 
+ bl[4] br[4] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_7 
+ bl[5] br[5] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_8 
+ bl[6] br[6] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_9 
+ bl[7] br[7] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_10 
+ bl[8] br[8] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_11 
+ bl[9] br[9] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_12 
+ bl[10] br[10] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_13 
+ bl[11] br[11] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_14 
+ bl[12] br[12] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_15 
+ bl[13] br[13] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_16 
+ bl[14] br[14] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_17 
+ bl[15] br[15] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_18 
+ bl[16] br[16] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_19 
+ bl[17] br[17] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_20 
+ bl[18] br[18] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_21 
+ bl[19] br[19] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_22 
+ bl[20] br[20] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_23 
+ bl[21] br[21] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_24 
+ bl[22] br[22] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_25 
+ bl[23] br[23] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_26 
+ bl[24] br[24] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_27 
+ bl[25] br[25] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_28 
+ bl[26] br[26] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_29 
+ bl[27] br[27] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_30 
+ bl[28] br[28] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_31 
+ bl[29] br[29] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_32 
+ bl[30] br[30] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_33 
+ bl[31] br[31] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_34 
+ bl[32] br[32] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_35 
+ bl[33] br[33] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_36 
+ bl[34] br[34] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_37 
+ bl[35] br[35] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_38 
+ bl[36] br[36] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_39 
+ bl[37] br[37] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_40 
+ bl[38] br[38] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_41 
+ bl[39] br[39] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_42 
+ bl[40] br[40] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_43 
+ bl[41] br[41] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_44 
+ bl[42] br[42] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_45 
+ bl[43] br[43] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_46 
+ bl[44] br[44] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_47 
+ bl[45] br[45] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_48 
+ bl[46] br[46] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_49 
+ bl[47] br[47] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_50 
+ bl[48] br[48] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_51 
+ bl[49] br[49] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_52 
+ bl[50] br[50] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_53 
+ bl[51] br[51] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_54 
+ bl[52] br[52] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_55 
+ bl[53] br[53] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_56 
+ bl[54] br[54] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_57 
+ bl[55] br[55] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_58 
+ bl[56] br[56] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_59 
+ bl[57] br[57] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_60 
+ bl[58] br[58] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_61 
+ bl[59] br[59] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_62 
+ bl[60] br[60] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_63 
+ bl[61] br[61] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_64 
+ bl[62] br[62] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_65 
+ bl[63] br[63] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_66 
+ bl[64] br[64] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_67 
+ bl[65] br[65] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_68 
+ bl[66] br[66] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_69 
+ bl[67] br[67] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_70 
+ bl[68] br[68] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_71 
+ bl[69] br[69] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_72 
+ bl[70] br[70] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_73 
+ bl[71] br[71] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_74 
+ bl[72] br[72] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_75 
+ bl[73] br[73] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_76 
+ bl[74] br[74] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_77 
+ bl[75] br[75] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_78 
+ bl[76] br[76] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_79 
+ bl[77] br[77] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_80 
+ bl[78] br[78] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_81 
+ bl[79] br[79] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_82 
+ bl[80] br[80] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_83 
+ bl[81] br[81] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_84 
+ bl[82] br[82] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_85 
+ bl[83] br[83] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_86 
+ bl[84] br[84] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_87 
+ bl[85] br[85] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_88 
+ bl[86] br[86] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_89 
+ bl[87] br[87] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_90 
+ bl[88] br[88] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_91 
+ bl[89] br[89] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_92 
+ bl[90] br[90] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_93 
+ bl[91] br[91] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_94 
+ bl[92] br[92] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_95 
+ bl[93] br[93] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_96 
+ bl[94] br[94] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_97 
+ bl[95] br[95] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_98 
+ bl[96] br[96] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_99 
+ bl[97] br[97] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_100 
+ bl[98] br[98] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_101 
+ bl[99] br[99] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_102 
+ bl[100] br[100] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_103 
+ bl[101] br[101] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_104 
+ bl[102] br[102] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_105 
+ bl[103] br[103] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_106 
+ bl[104] br[104] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_107 
+ bl[105] br[105] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_108 
+ bl[106] br[106] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_109 
+ bl[107] br[107] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_110 
+ bl[108] br[108] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_111 
+ bl[109] br[109] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_112 
+ bl[110] br[110] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_113 
+ bl[111] br[111] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_114 
+ bl[112] br[112] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_115 
+ bl[113] br[113] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_116 
+ bl[114] br[114] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_117 
+ bl[115] br[115] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_118 
+ bl[116] br[116] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_119 
+ bl[117] br[117] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_120 
+ bl[118] br[118] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_121 
+ bl[119] br[119] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_122 
+ bl[120] br[120] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_123 
+ bl[121] br[121] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_124 
+ bl[122] br[122] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_125 
+ bl[123] br[123] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_126 
+ bl[124] br[124] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_127 
+ bl[125] br[125] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_128 
+ bl[126] br[126] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_129 
+ bl[127] br[127] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_130 
+ vdd vdd vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_131 
+ vdd vdd vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_0 
+ vdd vdd vss vdd vpb vnb wl[58] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_60_1 
+ rbl rbr vss vdd vpb vnb wl[58] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_60_2 
+ bl[0] br[0] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_3 
+ bl[1] br[1] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_4 
+ bl[2] br[2] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_5 
+ bl[3] br[3] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_6 
+ bl[4] br[4] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_7 
+ bl[5] br[5] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_8 
+ bl[6] br[6] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_9 
+ bl[7] br[7] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_10 
+ bl[8] br[8] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_11 
+ bl[9] br[9] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_12 
+ bl[10] br[10] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_13 
+ bl[11] br[11] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_14 
+ bl[12] br[12] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_15 
+ bl[13] br[13] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_16 
+ bl[14] br[14] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_17 
+ bl[15] br[15] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_18 
+ bl[16] br[16] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_19 
+ bl[17] br[17] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_20 
+ bl[18] br[18] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_21 
+ bl[19] br[19] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_22 
+ bl[20] br[20] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_23 
+ bl[21] br[21] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_24 
+ bl[22] br[22] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_25 
+ bl[23] br[23] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_26 
+ bl[24] br[24] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_27 
+ bl[25] br[25] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_28 
+ bl[26] br[26] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_29 
+ bl[27] br[27] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_30 
+ bl[28] br[28] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_31 
+ bl[29] br[29] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_32 
+ bl[30] br[30] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_33 
+ bl[31] br[31] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_34 
+ bl[32] br[32] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_35 
+ bl[33] br[33] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_36 
+ bl[34] br[34] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_37 
+ bl[35] br[35] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_38 
+ bl[36] br[36] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_39 
+ bl[37] br[37] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_40 
+ bl[38] br[38] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_41 
+ bl[39] br[39] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_42 
+ bl[40] br[40] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_43 
+ bl[41] br[41] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_44 
+ bl[42] br[42] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_45 
+ bl[43] br[43] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_46 
+ bl[44] br[44] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_47 
+ bl[45] br[45] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_48 
+ bl[46] br[46] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_49 
+ bl[47] br[47] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_50 
+ bl[48] br[48] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_51 
+ bl[49] br[49] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_52 
+ bl[50] br[50] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_53 
+ bl[51] br[51] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_54 
+ bl[52] br[52] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_55 
+ bl[53] br[53] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_56 
+ bl[54] br[54] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_57 
+ bl[55] br[55] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_58 
+ bl[56] br[56] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_59 
+ bl[57] br[57] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_60 
+ bl[58] br[58] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_61 
+ bl[59] br[59] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_62 
+ bl[60] br[60] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_63 
+ bl[61] br[61] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_64 
+ bl[62] br[62] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_65 
+ bl[63] br[63] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_66 
+ bl[64] br[64] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_67 
+ bl[65] br[65] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_68 
+ bl[66] br[66] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_69 
+ bl[67] br[67] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_70 
+ bl[68] br[68] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_71 
+ bl[69] br[69] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_72 
+ bl[70] br[70] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_73 
+ bl[71] br[71] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_74 
+ bl[72] br[72] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_75 
+ bl[73] br[73] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_76 
+ bl[74] br[74] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_77 
+ bl[75] br[75] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_78 
+ bl[76] br[76] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_79 
+ bl[77] br[77] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_80 
+ bl[78] br[78] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_81 
+ bl[79] br[79] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_82 
+ bl[80] br[80] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_83 
+ bl[81] br[81] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_84 
+ bl[82] br[82] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_85 
+ bl[83] br[83] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_86 
+ bl[84] br[84] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_87 
+ bl[85] br[85] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_88 
+ bl[86] br[86] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_89 
+ bl[87] br[87] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_90 
+ bl[88] br[88] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_91 
+ bl[89] br[89] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_92 
+ bl[90] br[90] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_93 
+ bl[91] br[91] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_94 
+ bl[92] br[92] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_95 
+ bl[93] br[93] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_96 
+ bl[94] br[94] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_97 
+ bl[95] br[95] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_98 
+ bl[96] br[96] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_99 
+ bl[97] br[97] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_100 
+ bl[98] br[98] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_101 
+ bl[99] br[99] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_102 
+ bl[100] br[100] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_103 
+ bl[101] br[101] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_104 
+ bl[102] br[102] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_105 
+ bl[103] br[103] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_106 
+ bl[104] br[104] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_107 
+ bl[105] br[105] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_108 
+ bl[106] br[106] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_109 
+ bl[107] br[107] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_110 
+ bl[108] br[108] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_111 
+ bl[109] br[109] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_112 
+ bl[110] br[110] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_113 
+ bl[111] br[111] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_114 
+ bl[112] br[112] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_115 
+ bl[113] br[113] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_116 
+ bl[114] br[114] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_117 
+ bl[115] br[115] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_118 
+ bl[116] br[116] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_119 
+ bl[117] br[117] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_120 
+ bl[118] br[118] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_121 
+ bl[119] br[119] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_122 
+ bl[120] br[120] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_123 
+ bl[121] br[121] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_124 
+ bl[122] br[122] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_125 
+ bl[123] br[123] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_126 
+ bl[124] br[124] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_127 
+ bl[125] br[125] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_128 
+ bl[126] br[126] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_129 
+ bl[127] br[127] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_130 
+ vdd vdd vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_131 
+ vdd vdd vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_0 
+ vdd vdd vss vdd vpb vnb wl[59] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_61_1 
+ rbl rbr vss vdd vpb vnb wl[59] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_61_2 
+ bl[0] br[0] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_3 
+ bl[1] br[1] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_4 
+ bl[2] br[2] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_5 
+ bl[3] br[3] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_6 
+ bl[4] br[4] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_7 
+ bl[5] br[5] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_8 
+ bl[6] br[6] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_9 
+ bl[7] br[7] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_10 
+ bl[8] br[8] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_11 
+ bl[9] br[9] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_12 
+ bl[10] br[10] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_13 
+ bl[11] br[11] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_14 
+ bl[12] br[12] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_15 
+ bl[13] br[13] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_16 
+ bl[14] br[14] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_17 
+ bl[15] br[15] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_18 
+ bl[16] br[16] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_19 
+ bl[17] br[17] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_20 
+ bl[18] br[18] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_21 
+ bl[19] br[19] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_22 
+ bl[20] br[20] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_23 
+ bl[21] br[21] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_24 
+ bl[22] br[22] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_25 
+ bl[23] br[23] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_26 
+ bl[24] br[24] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_27 
+ bl[25] br[25] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_28 
+ bl[26] br[26] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_29 
+ bl[27] br[27] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_30 
+ bl[28] br[28] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_31 
+ bl[29] br[29] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_32 
+ bl[30] br[30] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_33 
+ bl[31] br[31] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_34 
+ bl[32] br[32] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_35 
+ bl[33] br[33] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_36 
+ bl[34] br[34] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_37 
+ bl[35] br[35] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_38 
+ bl[36] br[36] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_39 
+ bl[37] br[37] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_40 
+ bl[38] br[38] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_41 
+ bl[39] br[39] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_42 
+ bl[40] br[40] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_43 
+ bl[41] br[41] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_44 
+ bl[42] br[42] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_45 
+ bl[43] br[43] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_46 
+ bl[44] br[44] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_47 
+ bl[45] br[45] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_48 
+ bl[46] br[46] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_49 
+ bl[47] br[47] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_50 
+ bl[48] br[48] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_51 
+ bl[49] br[49] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_52 
+ bl[50] br[50] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_53 
+ bl[51] br[51] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_54 
+ bl[52] br[52] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_55 
+ bl[53] br[53] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_56 
+ bl[54] br[54] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_57 
+ bl[55] br[55] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_58 
+ bl[56] br[56] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_59 
+ bl[57] br[57] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_60 
+ bl[58] br[58] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_61 
+ bl[59] br[59] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_62 
+ bl[60] br[60] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_63 
+ bl[61] br[61] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_64 
+ bl[62] br[62] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_65 
+ bl[63] br[63] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_66 
+ bl[64] br[64] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_67 
+ bl[65] br[65] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_68 
+ bl[66] br[66] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_69 
+ bl[67] br[67] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_70 
+ bl[68] br[68] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_71 
+ bl[69] br[69] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_72 
+ bl[70] br[70] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_73 
+ bl[71] br[71] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_74 
+ bl[72] br[72] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_75 
+ bl[73] br[73] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_76 
+ bl[74] br[74] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_77 
+ bl[75] br[75] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_78 
+ bl[76] br[76] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_79 
+ bl[77] br[77] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_80 
+ bl[78] br[78] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_81 
+ bl[79] br[79] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_82 
+ bl[80] br[80] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_83 
+ bl[81] br[81] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_84 
+ bl[82] br[82] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_85 
+ bl[83] br[83] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_86 
+ bl[84] br[84] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_87 
+ bl[85] br[85] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_88 
+ bl[86] br[86] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_89 
+ bl[87] br[87] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_90 
+ bl[88] br[88] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_91 
+ bl[89] br[89] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_92 
+ bl[90] br[90] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_93 
+ bl[91] br[91] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_94 
+ bl[92] br[92] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_95 
+ bl[93] br[93] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_96 
+ bl[94] br[94] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_97 
+ bl[95] br[95] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_98 
+ bl[96] br[96] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_99 
+ bl[97] br[97] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_100 
+ bl[98] br[98] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_101 
+ bl[99] br[99] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_102 
+ bl[100] br[100] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_103 
+ bl[101] br[101] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_104 
+ bl[102] br[102] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_105 
+ bl[103] br[103] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_106 
+ bl[104] br[104] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_107 
+ bl[105] br[105] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_108 
+ bl[106] br[106] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_109 
+ bl[107] br[107] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_110 
+ bl[108] br[108] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_111 
+ bl[109] br[109] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_112 
+ bl[110] br[110] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_113 
+ bl[111] br[111] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_114 
+ bl[112] br[112] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_115 
+ bl[113] br[113] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_116 
+ bl[114] br[114] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_117 
+ bl[115] br[115] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_118 
+ bl[116] br[116] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_119 
+ bl[117] br[117] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_120 
+ bl[118] br[118] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_121 
+ bl[119] br[119] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_122 
+ bl[120] br[120] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_123 
+ bl[121] br[121] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_124 
+ bl[122] br[122] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_125 
+ bl[123] br[123] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_126 
+ bl[124] br[124] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_127 
+ bl[125] br[125] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_128 
+ bl[126] br[126] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_129 
+ bl[127] br[127] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_130 
+ vdd vdd vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_131 
+ vdd vdd vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_0 
+ vdd vdd vss vdd vpb vnb wl[60] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_62_1 
+ rbl rbr vss vdd vpb vnb wl[60] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_62_2 
+ bl[0] br[0] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_3 
+ bl[1] br[1] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_4 
+ bl[2] br[2] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_5 
+ bl[3] br[3] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_6 
+ bl[4] br[4] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_7 
+ bl[5] br[5] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_8 
+ bl[6] br[6] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_9 
+ bl[7] br[7] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_10 
+ bl[8] br[8] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_11 
+ bl[9] br[9] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_12 
+ bl[10] br[10] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_13 
+ bl[11] br[11] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_14 
+ bl[12] br[12] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_15 
+ bl[13] br[13] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_16 
+ bl[14] br[14] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_17 
+ bl[15] br[15] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_18 
+ bl[16] br[16] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_19 
+ bl[17] br[17] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_20 
+ bl[18] br[18] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_21 
+ bl[19] br[19] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_22 
+ bl[20] br[20] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_23 
+ bl[21] br[21] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_24 
+ bl[22] br[22] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_25 
+ bl[23] br[23] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_26 
+ bl[24] br[24] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_27 
+ bl[25] br[25] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_28 
+ bl[26] br[26] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_29 
+ bl[27] br[27] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_30 
+ bl[28] br[28] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_31 
+ bl[29] br[29] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_32 
+ bl[30] br[30] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_33 
+ bl[31] br[31] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_34 
+ bl[32] br[32] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_35 
+ bl[33] br[33] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_36 
+ bl[34] br[34] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_37 
+ bl[35] br[35] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_38 
+ bl[36] br[36] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_39 
+ bl[37] br[37] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_40 
+ bl[38] br[38] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_41 
+ bl[39] br[39] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_42 
+ bl[40] br[40] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_43 
+ bl[41] br[41] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_44 
+ bl[42] br[42] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_45 
+ bl[43] br[43] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_46 
+ bl[44] br[44] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_47 
+ bl[45] br[45] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_48 
+ bl[46] br[46] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_49 
+ bl[47] br[47] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_50 
+ bl[48] br[48] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_51 
+ bl[49] br[49] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_52 
+ bl[50] br[50] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_53 
+ bl[51] br[51] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_54 
+ bl[52] br[52] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_55 
+ bl[53] br[53] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_56 
+ bl[54] br[54] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_57 
+ bl[55] br[55] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_58 
+ bl[56] br[56] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_59 
+ bl[57] br[57] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_60 
+ bl[58] br[58] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_61 
+ bl[59] br[59] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_62 
+ bl[60] br[60] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_63 
+ bl[61] br[61] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_64 
+ bl[62] br[62] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_65 
+ bl[63] br[63] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_66 
+ bl[64] br[64] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_67 
+ bl[65] br[65] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_68 
+ bl[66] br[66] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_69 
+ bl[67] br[67] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_70 
+ bl[68] br[68] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_71 
+ bl[69] br[69] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_72 
+ bl[70] br[70] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_73 
+ bl[71] br[71] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_74 
+ bl[72] br[72] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_75 
+ bl[73] br[73] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_76 
+ bl[74] br[74] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_77 
+ bl[75] br[75] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_78 
+ bl[76] br[76] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_79 
+ bl[77] br[77] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_80 
+ bl[78] br[78] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_81 
+ bl[79] br[79] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_82 
+ bl[80] br[80] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_83 
+ bl[81] br[81] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_84 
+ bl[82] br[82] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_85 
+ bl[83] br[83] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_86 
+ bl[84] br[84] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_87 
+ bl[85] br[85] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_88 
+ bl[86] br[86] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_89 
+ bl[87] br[87] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_90 
+ bl[88] br[88] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_91 
+ bl[89] br[89] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_92 
+ bl[90] br[90] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_93 
+ bl[91] br[91] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_94 
+ bl[92] br[92] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_95 
+ bl[93] br[93] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_96 
+ bl[94] br[94] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_97 
+ bl[95] br[95] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_98 
+ bl[96] br[96] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_99 
+ bl[97] br[97] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_100 
+ bl[98] br[98] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_101 
+ bl[99] br[99] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_102 
+ bl[100] br[100] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_103 
+ bl[101] br[101] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_104 
+ bl[102] br[102] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_105 
+ bl[103] br[103] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_106 
+ bl[104] br[104] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_107 
+ bl[105] br[105] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_108 
+ bl[106] br[106] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_109 
+ bl[107] br[107] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_110 
+ bl[108] br[108] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_111 
+ bl[109] br[109] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_112 
+ bl[110] br[110] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_113 
+ bl[111] br[111] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_114 
+ bl[112] br[112] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_115 
+ bl[113] br[113] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_116 
+ bl[114] br[114] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_117 
+ bl[115] br[115] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_118 
+ bl[116] br[116] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_119 
+ bl[117] br[117] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_120 
+ bl[118] br[118] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_121 
+ bl[119] br[119] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_122 
+ bl[120] br[120] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_123 
+ bl[121] br[121] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_124 
+ bl[122] br[122] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_125 
+ bl[123] br[123] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_126 
+ bl[124] br[124] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_127 
+ bl[125] br[125] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_128 
+ bl[126] br[126] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_129 
+ bl[127] br[127] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_130 
+ vdd vdd vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_131 
+ vdd vdd vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_0 
+ vdd vdd vss vdd vpb vnb wl[61] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_63_1 
+ rbl rbr vss vdd vpb vnb wl[61] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_63_2 
+ bl[0] br[0] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_3 
+ bl[1] br[1] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_4 
+ bl[2] br[2] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_5 
+ bl[3] br[3] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_6 
+ bl[4] br[4] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_7 
+ bl[5] br[5] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_8 
+ bl[6] br[6] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_9 
+ bl[7] br[7] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_10 
+ bl[8] br[8] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_11 
+ bl[9] br[9] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_12 
+ bl[10] br[10] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_13 
+ bl[11] br[11] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_14 
+ bl[12] br[12] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_15 
+ bl[13] br[13] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_16 
+ bl[14] br[14] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_17 
+ bl[15] br[15] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_18 
+ bl[16] br[16] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_19 
+ bl[17] br[17] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_20 
+ bl[18] br[18] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_21 
+ bl[19] br[19] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_22 
+ bl[20] br[20] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_23 
+ bl[21] br[21] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_24 
+ bl[22] br[22] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_25 
+ bl[23] br[23] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_26 
+ bl[24] br[24] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_27 
+ bl[25] br[25] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_28 
+ bl[26] br[26] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_29 
+ bl[27] br[27] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_30 
+ bl[28] br[28] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_31 
+ bl[29] br[29] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_32 
+ bl[30] br[30] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_33 
+ bl[31] br[31] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_34 
+ bl[32] br[32] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_35 
+ bl[33] br[33] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_36 
+ bl[34] br[34] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_37 
+ bl[35] br[35] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_38 
+ bl[36] br[36] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_39 
+ bl[37] br[37] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_40 
+ bl[38] br[38] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_41 
+ bl[39] br[39] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_42 
+ bl[40] br[40] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_43 
+ bl[41] br[41] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_44 
+ bl[42] br[42] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_45 
+ bl[43] br[43] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_46 
+ bl[44] br[44] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_47 
+ bl[45] br[45] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_48 
+ bl[46] br[46] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_49 
+ bl[47] br[47] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_50 
+ bl[48] br[48] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_51 
+ bl[49] br[49] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_52 
+ bl[50] br[50] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_53 
+ bl[51] br[51] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_54 
+ bl[52] br[52] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_55 
+ bl[53] br[53] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_56 
+ bl[54] br[54] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_57 
+ bl[55] br[55] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_58 
+ bl[56] br[56] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_59 
+ bl[57] br[57] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_60 
+ bl[58] br[58] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_61 
+ bl[59] br[59] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_62 
+ bl[60] br[60] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_63 
+ bl[61] br[61] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_64 
+ bl[62] br[62] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_65 
+ bl[63] br[63] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_66 
+ bl[64] br[64] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_67 
+ bl[65] br[65] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_68 
+ bl[66] br[66] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_69 
+ bl[67] br[67] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_70 
+ bl[68] br[68] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_71 
+ bl[69] br[69] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_72 
+ bl[70] br[70] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_73 
+ bl[71] br[71] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_74 
+ bl[72] br[72] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_75 
+ bl[73] br[73] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_76 
+ bl[74] br[74] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_77 
+ bl[75] br[75] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_78 
+ bl[76] br[76] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_79 
+ bl[77] br[77] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_80 
+ bl[78] br[78] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_81 
+ bl[79] br[79] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_82 
+ bl[80] br[80] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_83 
+ bl[81] br[81] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_84 
+ bl[82] br[82] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_85 
+ bl[83] br[83] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_86 
+ bl[84] br[84] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_87 
+ bl[85] br[85] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_88 
+ bl[86] br[86] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_89 
+ bl[87] br[87] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_90 
+ bl[88] br[88] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_91 
+ bl[89] br[89] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_92 
+ bl[90] br[90] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_93 
+ bl[91] br[91] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_94 
+ bl[92] br[92] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_95 
+ bl[93] br[93] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_96 
+ bl[94] br[94] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_97 
+ bl[95] br[95] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_98 
+ bl[96] br[96] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_99 
+ bl[97] br[97] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_100 
+ bl[98] br[98] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_101 
+ bl[99] br[99] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_102 
+ bl[100] br[100] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_103 
+ bl[101] br[101] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_104 
+ bl[102] br[102] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_105 
+ bl[103] br[103] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_106 
+ bl[104] br[104] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_107 
+ bl[105] br[105] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_108 
+ bl[106] br[106] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_109 
+ bl[107] br[107] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_110 
+ bl[108] br[108] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_111 
+ bl[109] br[109] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_112 
+ bl[110] br[110] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_113 
+ bl[111] br[111] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_114 
+ bl[112] br[112] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_115 
+ bl[113] br[113] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_116 
+ bl[114] br[114] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_117 
+ bl[115] br[115] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_118 
+ bl[116] br[116] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_119 
+ bl[117] br[117] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_120 
+ bl[118] br[118] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_121 
+ bl[119] br[119] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_122 
+ bl[120] br[120] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_123 
+ bl[121] br[121] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_124 
+ bl[122] br[122] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_125 
+ bl[123] br[123] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_126 
+ bl[124] br[124] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_127 
+ bl[125] br[125] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_128 
+ bl[126] br[126] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_129 
+ bl[127] br[127] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_130 
+ vdd vdd vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_131 
+ vdd vdd vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_0 
+ vdd vdd vss vdd vpb vnb wl[62] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_64_1 
+ rbl rbr vss vdd vpb vnb wl[62] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_64_2 
+ bl[0] br[0] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_3 
+ bl[1] br[1] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_4 
+ bl[2] br[2] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_5 
+ bl[3] br[3] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_6 
+ bl[4] br[4] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_7 
+ bl[5] br[5] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_8 
+ bl[6] br[6] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_9 
+ bl[7] br[7] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_10 
+ bl[8] br[8] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_11 
+ bl[9] br[9] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_12 
+ bl[10] br[10] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_13 
+ bl[11] br[11] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_14 
+ bl[12] br[12] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_15 
+ bl[13] br[13] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_16 
+ bl[14] br[14] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_17 
+ bl[15] br[15] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_18 
+ bl[16] br[16] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_19 
+ bl[17] br[17] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_20 
+ bl[18] br[18] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_21 
+ bl[19] br[19] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_22 
+ bl[20] br[20] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_23 
+ bl[21] br[21] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_24 
+ bl[22] br[22] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_25 
+ bl[23] br[23] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_26 
+ bl[24] br[24] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_27 
+ bl[25] br[25] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_28 
+ bl[26] br[26] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_29 
+ bl[27] br[27] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_30 
+ bl[28] br[28] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_31 
+ bl[29] br[29] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_32 
+ bl[30] br[30] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_33 
+ bl[31] br[31] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_34 
+ bl[32] br[32] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_35 
+ bl[33] br[33] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_36 
+ bl[34] br[34] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_37 
+ bl[35] br[35] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_38 
+ bl[36] br[36] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_39 
+ bl[37] br[37] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_40 
+ bl[38] br[38] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_41 
+ bl[39] br[39] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_42 
+ bl[40] br[40] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_43 
+ bl[41] br[41] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_44 
+ bl[42] br[42] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_45 
+ bl[43] br[43] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_46 
+ bl[44] br[44] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_47 
+ bl[45] br[45] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_48 
+ bl[46] br[46] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_49 
+ bl[47] br[47] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_50 
+ bl[48] br[48] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_51 
+ bl[49] br[49] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_52 
+ bl[50] br[50] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_53 
+ bl[51] br[51] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_54 
+ bl[52] br[52] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_55 
+ bl[53] br[53] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_56 
+ bl[54] br[54] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_57 
+ bl[55] br[55] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_58 
+ bl[56] br[56] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_59 
+ bl[57] br[57] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_60 
+ bl[58] br[58] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_61 
+ bl[59] br[59] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_62 
+ bl[60] br[60] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_63 
+ bl[61] br[61] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_64 
+ bl[62] br[62] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_65 
+ bl[63] br[63] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_66 
+ bl[64] br[64] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_67 
+ bl[65] br[65] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_68 
+ bl[66] br[66] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_69 
+ bl[67] br[67] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_70 
+ bl[68] br[68] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_71 
+ bl[69] br[69] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_72 
+ bl[70] br[70] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_73 
+ bl[71] br[71] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_74 
+ bl[72] br[72] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_75 
+ bl[73] br[73] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_76 
+ bl[74] br[74] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_77 
+ bl[75] br[75] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_78 
+ bl[76] br[76] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_79 
+ bl[77] br[77] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_80 
+ bl[78] br[78] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_81 
+ bl[79] br[79] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_82 
+ bl[80] br[80] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_83 
+ bl[81] br[81] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_84 
+ bl[82] br[82] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_85 
+ bl[83] br[83] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_86 
+ bl[84] br[84] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_87 
+ bl[85] br[85] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_88 
+ bl[86] br[86] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_89 
+ bl[87] br[87] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_90 
+ bl[88] br[88] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_91 
+ bl[89] br[89] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_92 
+ bl[90] br[90] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_93 
+ bl[91] br[91] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_94 
+ bl[92] br[92] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_95 
+ bl[93] br[93] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_96 
+ bl[94] br[94] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_97 
+ bl[95] br[95] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_98 
+ bl[96] br[96] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_99 
+ bl[97] br[97] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_100 
+ bl[98] br[98] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_101 
+ bl[99] br[99] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_102 
+ bl[100] br[100] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_103 
+ bl[101] br[101] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_104 
+ bl[102] br[102] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_105 
+ bl[103] br[103] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_106 
+ bl[104] br[104] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_107 
+ bl[105] br[105] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_108 
+ bl[106] br[106] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_109 
+ bl[107] br[107] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_110 
+ bl[108] br[108] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_111 
+ bl[109] br[109] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_112 
+ bl[110] br[110] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_113 
+ bl[111] br[111] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_114 
+ bl[112] br[112] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_115 
+ bl[113] br[113] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_116 
+ bl[114] br[114] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_117 
+ bl[115] br[115] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_118 
+ bl[116] br[116] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_119 
+ bl[117] br[117] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_120 
+ bl[118] br[118] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_121 
+ bl[119] br[119] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_122 
+ bl[120] br[120] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_123 
+ bl[121] br[121] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_124 
+ bl[122] br[122] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_125 
+ bl[123] br[123] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_126 
+ bl[124] br[124] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_127 
+ bl[125] br[125] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_128 
+ bl[126] br[126] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_129 
+ bl[127] br[127] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_130 
+ vdd vdd vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_131 
+ vdd vdd vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_0 
+ vdd vdd vss vdd vpb vnb wl[63] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_65_1 
+ rbl rbr vss vdd vpb vnb wl[63] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_65_2 
+ bl[0] br[0] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_3 
+ bl[1] br[1] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_4 
+ bl[2] br[2] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_5 
+ bl[3] br[3] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_6 
+ bl[4] br[4] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_7 
+ bl[5] br[5] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_8 
+ bl[6] br[6] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_9 
+ bl[7] br[7] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_10 
+ bl[8] br[8] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_11 
+ bl[9] br[9] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_12 
+ bl[10] br[10] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_13 
+ bl[11] br[11] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_14 
+ bl[12] br[12] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_15 
+ bl[13] br[13] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_16 
+ bl[14] br[14] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_17 
+ bl[15] br[15] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_18 
+ bl[16] br[16] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_19 
+ bl[17] br[17] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_20 
+ bl[18] br[18] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_21 
+ bl[19] br[19] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_22 
+ bl[20] br[20] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_23 
+ bl[21] br[21] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_24 
+ bl[22] br[22] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_25 
+ bl[23] br[23] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_26 
+ bl[24] br[24] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_27 
+ bl[25] br[25] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_28 
+ bl[26] br[26] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_29 
+ bl[27] br[27] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_30 
+ bl[28] br[28] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_31 
+ bl[29] br[29] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_32 
+ bl[30] br[30] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_33 
+ bl[31] br[31] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_34 
+ bl[32] br[32] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_35 
+ bl[33] br[33] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_36 
+ bl[34] br[34] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_37 
+ bl[35] br[35] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_38 
+ bl[36] br[36] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_39 
+ bl[37] br[37] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_40 
+ bl[38] br[38] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_41 
+ bl[39] br[39] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_42 
+ bl[40] br[40] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_43 
+ bl[41] br[41] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_44 
+ bl[42] br[42] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_45 
+ bl[43] br[43] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_46 
+ bl[44] br[44] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_47 
+ bl[45] br[45] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_48 
+ bl[46] br[46] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_49 
+ bl[47] br[47] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_50 
+ bl[48] br[48] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_51 
+ bl[49] br[49] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_52 
+ bl[50] br[50] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_53 
+ bl[51] br[51] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_54 
+ bl[52] br[52] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_55 
+ bl[53] br[53] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_56 
+ bl[54] br[54] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_57 
+ bl[55] br[55] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_58 
+ bl[56] br[56] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_59 
+ bl[57] br[57] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_60 
+ bl[58] br[58] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_61 
+ bl[59] br[59] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_62 
+ bl[60] br[60] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_63 
+ bl[61] br[61] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_64 
+ bl[62] br[62] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_65 
+ bl[63] br[63] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_66 
+ bl[64] br[64] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_67 
+ bl[65] br[65] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_68 
+ bl[66] br[66] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_69 
+ bl[67] br[67] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_70 
+ bl[68] br[68] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_71 
+ bl[69] br[69] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_72 
+ bl[70] br[70] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_73 
+ bl[71] br[71] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_74 
+ bl[72] br[72] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_75 
+ bl[73] br[73] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_76 
+ bl[74] br[74] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_77 
+ bl[75] br[75] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_78 
+ bl[76] br[76] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_79 
+ bl[77] br[77] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_80 
+ bl[78] br[78] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_81 
+ bl[79] br[79] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_82 
+ bl[80] br[80] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_83 
+ bl[81] br[81] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_84 
+ bl[82] br[82] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_85 
+ bl[83] br[83] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_86 
+ bl[84] br[84] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_87 
+ bl[85] br[85] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_88 
+ bl[86] br[86] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_89 
+ bl[87] br[87] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_90 
+ bl[88] br[88] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_91 
+ bl[89] br[89] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_92 
+ bl[90] br[90] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_93 
+ bl[91] br[91] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_94 
+ bl[92] br[92] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_95 
+ bl[93] br[93] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_96 
+ bl[94] br[94] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_97 
+ bl[95] br[95] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_98 
+ bl[96] br[96] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_99 
+ bl[97] br[97] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_100 
+ bl[98] br[98] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_101 
+ bl[99] br[99] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_102 
+ bl[100] br[100] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_103 
+ bl[101] br[101] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_104 
+ bl[102] br[102] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_105 
+ bl[103] br[103] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_106 
+ bl[104] br[104] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_107 
+ bl[105] br[105] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_108 
+ bl[106] br[106] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_109 
+ bl[107] br[107] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_110 
+ bl[108] br[108] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_111 
+ bl[109] br[109] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_112 
+ bl[110] br[110] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_113 
+ bl[111] br[111] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_114 
+ bl[112] br[112] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_115 
+ bl[113] br[113] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_116 
+ bl[114] br[114] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_117 
+ bl[115] br[115] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_118 
+ bl[116] br[116] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_119 
+ bl[117] br[117] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_120 
+ bl[118] br[118] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_121 
+ bl[119] br[119] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_122 
+ bl[120] br[120] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_123 
+ bl[121] br[121] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_124 
+ bl[122] br[122] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_125 
+ bl[123] br[123] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_126 
+ bl[124] br[124] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_127 
+ bl[125] br[125] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_128 
+ bl[126] br[126] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_129 
+ bl[127] br[127] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_130 
+ vdd vdd vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_131 
+ vdd vdd vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_130 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_131 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_130 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_131 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xcolend_0_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_0_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_bot 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_top 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_bot 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_top 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_bot 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_top 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_bot 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_top 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_bot 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_top 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_bot 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_top 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_bot 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_top 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_bot 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_top 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_bot 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_top 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_bot 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_top 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_bot 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_top 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_bot 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_top 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_bot 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_top 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_bot 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_top 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_bot 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_top 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_bot 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_top 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_bot 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_top 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_bot 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_top 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_bot 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_top 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_bot 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_top 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_bot 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_top 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_bot 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_top 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_bot 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_top 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_bot 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_top 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_bot 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_top 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_bot 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_top 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_bot 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_top 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_bot 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_top 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_bot 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_top 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_bot 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_top 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_bot 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_top 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_bot 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_top 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_bot 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_top 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_bot 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_top 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_bot 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_top 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_bot 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_top 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_bot 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_top 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_bot 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_top 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_bot 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_top 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_bot 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_top 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_bot 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_top 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_bot 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_top 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_bot 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_top 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_bot 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_top 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_bot 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_top 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_bot 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_top 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_bot 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_top 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_bot 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_top 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_bot 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_top 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_bot 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_top 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_bot 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_top 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_bot 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_top 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_bot 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_top 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_bot 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_top 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_bot 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_top 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_bot 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_top 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_bot 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_top 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_bot 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_top 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_bot 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_top 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_bot 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_top 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_bot 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_top 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_bot 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_top 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_bot 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_top 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_bot 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_top 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_bot 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_top 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_bot 
+ br[64] vdd vss bl[64] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_top 
+ br[64] vdd vss bl[64] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_bot 
+ br[65] vdd vss bl[65] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_top 
+ br[65] vdd vss bl[65] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_68_bot 
+ br[66] vdd vss bl[66] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_68_top 
+ br[66] vdd vss bl[66] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_69_bot 
+ br[67] vdd vss bl[67] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_69_top 
+ br[67] vdd vss bl[67] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_70_bot 
+ br[68] vdd vss bl[68] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_70_top 
+ br[68] vdd vss bl[68] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_71_bot 
+ br[69] vdd vss bl[69] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_71_top 
+ br[69] vdd vss bl[69] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_72_bot 
+ br[70] vdd vss bl[70] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_72_top 
+ br[70] vdd vss bl[70] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_73_bot 
+ br[71] vdd vss bl[71] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_73_top 
+ br[71] vdd vss bl[71] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_74_bot 
+ br[72] vdd vss bl[72] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_74_top 
+ br[72] vdd vss bl[72] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_75_bot 
+ br[73] vdd vss bl[73] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_75_top 
+ br[73] vdd vss bl[73] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_76_bot 
+ br[74] vdd vss bl[74] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_76_top 
+ br[74] vdd vss bl[74] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_77_bot 
+ br[75] vdd vss bl[75] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_77_top 
+ br[75] vdd vss bl[75] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_78_bot 
+ br[76] vdd vss bl[76] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_78_top 
+ br[76] vdd vss bl[76] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_79_bot 
+ br[77] vdd vss bl[77] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_79_top 
+ br[77] vdd vss bl[77] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_80_bot 
+ br[78] vdd vss bl[78] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_80_top 
+ br[78] vdd vss bl[78] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_81_bot 
+ br[79] vdd vss bl[79] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_81_top 
+ br[79] vdd vss bl[79] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_82_bot 
+ br[80] vdd vss bl[80] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_82_top 
+ br[80] vdd vss bl[80] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_83_bot 
+ br[81] vdd vss bl[81] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_83_top 
+ br[81] vdd vss bl[81] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_84_bot 
+ br[82] vdd vss bl[82] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_84_top 
+ br[82] vdd vss bl[82] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_85_bot 
+ br[83] vdd vss bl[83] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_85_top 
+ br[83] vdd vss bl[83] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_86_bot 
+ br[84] vdd vss bl[84] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_86_top 
+ br[84] vdd vss bl[84] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_87_bot 
+ br[85] vdd vss bl[85] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_87_top 
+ br[85] vdd vss bl[85] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_88_bot 
+ br[86] vdd vss bl[86] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_88_top 
+ br[86] vdd vss bl[86] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_89_bot 
+ br[87] vdd vss bl[87] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_89_top 
+ br[87] vdd vss bl[87] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_90_bot 
+ br[88] vdd vss bl[88] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_90_top 
+ br[88] vdd vss bl[88] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_91_bot 
+ br[89] vdd vss bl[89] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_91_top 
+ br[89] vdd vss bl[89] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_92_bot 
+ br[90] vdd vss bl[90] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_92_top 
+ br[90] vdd vss bl[90] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_93_bot 
+ br[91] vdd vss bl[91] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_93_top 
+ br[91] vdd vss bl[91] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_94_bot 
+ br[92] vdd vss bl[92] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_94_top 
+ br[92] vdd vss bl[92] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_95_bot 
+ br[93] vdd vss bl[93] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_95_top 
+ br[93] vdd vss bl[93] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_96_bot 
+ br[94] vdd vss bl[94] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_96_top 
+ br[94] vdd vss bl[94] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_97_bot 
+ br[95] vdd vss bl[95] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_97_top 
+ br[95] vdd vss bl[95] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_98_bot 
+ br[96] vdd vss bl[96] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_98_top 
+ br[96] vdd vss bl[96] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_99_bot 
+ br[97] vdd vss bl[97] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_99_top 
+ br[97] vdd vss bl[97] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_100_bot 
+ br[98] vdd vss bl[98] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_100_top 
+ br[98] vdd vss bl[98] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_101_bot 
+ br[99] vdd vss bl[99] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_101_top 
+ br[99] vdd vss bl[99] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_102_bot 
+ br[100] vdd vss bl[100] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_102_top 
+ br[100] vdd vss bl[100] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_103_bot 
+ br[101] vdd vss bl[101] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_103_top 
+ br[101] vdd vss bl[101] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_104_bot 
+ br[102] vdd vss bl[102] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_104_top 
+ br[102] vdd vss bl[102] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_105_bot 
+ br[103] vdd vss bl[103] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_105_top 
+ br[103] vdd vss bl[103] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_106_bot 
+ br[104] vdd vss bl[104] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_106_top 
+ br[104] vdd vss bl[104] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_107_bot 
+ br[105] vdd vss bl[105] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_107_top 
+ br[105] vdd vss bl[105] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_108_bot 
+ br[106] vdd vss bl[106] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_108_top 
+ br[106] vdd vss bl[106] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_109_bot 
+ br[107] vdd vss bl[107] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_109_top 
+ br[107] vdd vss bl[107] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_110_bot 
+ br[108] vdd vss bl[108] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_110_top 
+ br[108] vdd vss bl[108] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_111_bot 
+ br[109] vdd vss bl[109] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_111_top 
+ br[109] vdd vss bl[109] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_112_bot 
+ br[110] vdd vss bl[110] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_112_top 
+ br[110] vdd vss bl[110] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_113_bot 
+ br[111] vdd vss bl[111] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_113_top 
+ br[111] vdd vss bl[111] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_114_bot 
+ br[112] vdd vss bl[112] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_114_top 
+ br[112] vdd vss bl[112] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_115_bot 
+ br[113] vdd vss bl[113] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_115_top 
+ br[113] vdd vss bl[113] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_116_bot 
+ br[114] vdd vss bl[114] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_116_top 
+ br[114] vdd vss bl[114] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_117_bot 
+ br[115] vdd vss bl[115] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_117_top 
+ br[115] vdd vss bl[115] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_118_bot 
+ br[116] vdd vss bl[116] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_118_top 
+ br[116] vdd vss bl[116] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_119_bot 
+ br[117] vdd vss bl[117] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_119_top 
+ br[117] vdd vss bl[117] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_120_bot 
+ br[118] vdd vss bl[118] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_120_top 
+ br[118] vdd vss bl[118] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_121_bot 
+ br[119] vdd vss bl[119] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_121_top 
+ br[119] vdd vss bl[119] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_122_bot 
+ br[120] vdd vss bl[120] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_122_top 
+ br[120] vdd vss bl[120] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_123_bot 
+ br[121] vdd vss bl[121] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_123_top 
+ br[121] vdd vss bl[121] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_124_bot 
+ br[122] vdd vss bl[122] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_124_top 
+ br[122] vdd vss bl[122] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_125_bot 
+ br[123] vdd vss bl[123] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_125_top 
+ br[123] vdd vss bl[123] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_126_bot 
+ br[124] vdd vss bl[124] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_126_top 
+ br[124] vdd vss bl[124] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_127_bot 
+ br[125] vdd vss bl[125] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_127_top 
+ br[125] vdd vss bl[125] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_128_bot 
+ br[126] vdd vss bl[126] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_128_top 
+ br[126] vdd vss bl[126] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_129_bot 
+ br[127] vdd vss bl[127] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_129_top 
+ br[127] vdd vss bl[127] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_130_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_130_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_131_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_131_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

.ENDS

.SUBCKT precharge 
+ vdd bl br en_b 

xbl_pull_up 
+ bl en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xbr_pull_up 
+ br en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xequalizer 
+ bl en_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

.ENDS

.SUBCKT precharge_array 
+ vdd en_b bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] 

xprecharge_0 
+ vdd bl[0] br[0] en_b 
+ precharge 
* No parameters

xprecharge_1 
+ vdd bl[1] br[1] en_b 
+ precharge 
* No parameters

xprecharge_2 
+ vdd bl[2] br[2] en_b 
+ precharge 
* No parameters

xprecharge_3 
+ vdd bl[3] br[3] en_b 
+ precharge 
* No parameters

xprecharge_4 
+ vdd bl[4] br[4] en_b 
+ precharge 
* No parameters

xprecharge_5 
+ vdd bl[5] br[5] en_b 
+ precharge 
* No parameters

xprecharge_6 
+ vdd bl[6] br[6] en_b 
+ precharge 
* No parameters

xprecharge_7 
+ vdd bl[7] br[7] en_b 
+ precharge 
* No parameters

xprecharge_8 
+ vdd bl[8] br[8] en_b 
+ precharge 
* No parameters

xprecharge_9 
+ vdd bl[9] br[9] en_b 
+ precharge 
* No parameters

xprecharge_10 
+ vdd bl[10] br[10] en_b 
+ precharge 
* No parameters

xprecharge_11 
+ vdd bl[11] br[11] en_b 
+ precharge 
* No parameters

xprecharge_12 
+ vdd bl[12] br[12] en_b 
+ precharge 
* No parameters

xprecharge_13 
+ vdd bl[13] br[13] en_b 
+ precharge 
* No parameters

xprecharge_14 
+ vdd bl[14] br[14] en_b 
+ precharge 
* No parameters

xprecharge_15 
+ vdd bl[15] br[15] en_b 
+ precharge 
* No parameters

xprecharge_16 
+ vdd bl[16] br[16] en_b 
+ precharge 
* No parameters

xprecharge_17 
+ vdd bl[17] br[17] en_b 
+ precharge 
* No parameters

xprecharge_18 
+ vdd bl[18] br[18] en_b 
+ precharge 
* No parameters

xprecharge_19 
+ vdd bl[19] br[19] en_b 
+ precharge 
* No parameters

xprecharge_20 
+ vdd bl[20] br[20] en_b 
+ precharge 
* No parameters

xprecharge_21 
+ vdd bl[21] br[21] en_b 
+ precharge 
* No parameters

xprecharge_22 
+ vdd bl[22] br[22] en_b 
+ precharge 
* No parameters

xprecharge_23 
+ vdd bl[23] br[23] en_b 
+ precharge 
* No parameters

xprecharge_24 
+ vdd bl[24] br[24] en_b 
+ precharge 
* No parameters

xprecharge_25 
+ vdd bl[25] br[25] en_b 
+ precharge 
* No parameters

xprecharge_26 
+ vdd bl[26] br[26] en_b 
+ precharge 
* No parameters

xprecharge_27 
+ vdd bl[27] br[27] en_b 
+ precharge 
* No parameters

xprecharge_28 
+ vdd bl[28] br[28] en_b 
+ precharge 
* No parameters

xprecharge_29 
+ vdd bl[29] br[29] en_b 
+ precharge 
* No parameters

xprecharge_30 
+ vdd bl[30] br[30] en_b 
+ precharge 
* No parameters

xprecharge_31 
+ vdd bl[31] br[31] en_b 
+ precharge 
* No parameters

xprecharge_32 
+ vdd bl[32] br[32] en_b 
+ precharge 
* No parameters

xprecharge_33 
+ vdd bl[33] br[33] en_b 
+ precharge 
* No parameters

xprecharge_34 
+ vdd bl[34] br[34] en_b 
+ precharge 
* No parameters

xprecharge_35 
+ vdd bl[35] br[35] en_b 
+ precharge 
* No parameters

xprecharge_36 
+ vdd bl[36] br[36] en_b 
+ precharge 
* No parameters

xprecharge_37 
+ vdd bl[37] br[37] en_b 
+ precharge 
* No parameters

xprecharge_38 
+ vdd bl[38] br[38] en_b 
+ precharge 
* No parameters

xprecharge_39 
+ vdd bl[39] br[39] en_b 
+ precharge 
* No parameters

xprecharge_40 
+ vdd bl[40] br[40] en_b 
+ precharge 
* No parameters

xprecharge_41 
+ vdd bl[41] br[41] en_b 
+ precharge 
* No parameters

xprecharge_42 
+ vdd bl[42] br[42] en_b 
+ precharge 
* No parameters

xprecharge_43 
+ vdd bl[43] br[43] en_b 
+ precharge 
* No parameters

xprecharge_44 
+ vdd bl[44] br[44] en_b 
+ precharge 
* No parameters

xprecharge_45 
+ vdd bl[45] br[45] en_b 
+ precharge 
* No parameters

xprecharge_46 
+ vdd bl[46] br[46] en_b 
+ precharge 
* No parameters

xprecharge_47 
+ vdd bl[47] br[47] en_b 
+ precharge 
* No parameters

xprecharge_48 
+ vdd bl[48] br[48] en_b 
+ precharge 
* No parameters

xprecharge_49 
+ vdd bl[49] br[49] en_b 
+ precharge 
* No parameters

xprecharge_50 
+ vdd bl[50] br[50] en_b 
+ precharge 
* No parameters

xprecharge_51 
+ vdd bl[51] br[51] en_b 
+ precharge 
* No parameters

xprecharge_52 
+ vdd bl[52] br[52] en_b 
+ precharge 
* No parameters

xprecharge_53 
+ vdd bl[53] br[53] en_b 
+ precharge 
* No parameters

xprecharge_54 
+ vdd bl[54] br[54] en_b 
+ precharge 
* No parameters

xprecharge_55 
+ vdd bl[55] br[55] en_b 
+ precharge 
* No parameters

xprecharge_56 
+ vdd bl[56] br[56] en_b 
+ precharge 
* No parameters

xprecharge_57 
+ vdd bl[57] br[57] en_b 
+ precharge 
* No parameters

xprecharge_58 
+ vdd bl[58] br[58] en_b 
+ precharge 
* No parameters

xprecharge_59 
+ vdd bl[59] br[59] en_b 
+ precharge 
* No parameters

xprecharge_60 
+ vdd bl[60] br[60] en_b 
+ precharge 
* No parameters

xprecharge_61 
+ vdd bl[61] br[61] en_b 
+ precharge 
* No parameters

xprecharge_62 
+ vdd bl[62] br[62] en_b 
+ precharge 
* No parameters

xprecharge_63 
+ vdd bl[63] br[63] en_b 
+ precharge 
* No parameters

xprecharge_64 
+ vdd bl[64] br[64] en_b 
+ precharge 
* No parameters

xprecharge_65 
+ vdd bl[65] br[65] en_b 
+ precharge 
* No parameters

xprecharge_66 
+ vdd bl[66] br[66] en_b 
+ precharge 
* No parameters

xprecharge_67 
+ vdd bl[67] br[67] en_b 
+ precharge 
* No parameters

xprecharge_68 
+ vdd bl[68] br[68] en_b 
+ precharge 
* No parameters

xprecharge_69 
+ vdd bl[69] br[69] en_b 
+ precharge 
* No parameters

xprecharge_70 
+ vdd bl[70] br[70] en_b 
+ precharge 
* No parameters

xprecharge_71 
+ vdd bl[71] br[71] en_b 
+ precharge 
* No parameters

xprecharge_72 
+ vdd bl[72] br[72] en_b 
+ precharge 
* No parameters

xprecharge_73 
+ vdd bl[73] br[73] en_b 
+ precharge 
* No parameters

xprecharge_74 
+ vdd bl[74] br[74] en_b 
+ precharge 
* No parameters

xprecharge_75 
+ vdd bl[75] br[75] en_b 
+ precharge 
* No parameters

xprecharge_76 
+ vdd bl[76] br[76] en_b 
+ precharge 
* No parameters

xprecharge_77 
+ vdd bl[77] br[77] en_b 
+ precharge 
* No parameters

xprecharge_78 
+ vdd bl[78] br[78] en_b 
+ precharge 
* No parameters

xprecharge_79 
+ vdd bl[79] br[79] en_b 
+ precharge 
* No parameters

xprecharge_80 
+ vdd bl[80] br[80] en_b 
+ precharge 
* No parameters

xprecharge_81 
+ vdd bl[81] br[81] en_b 
+ precharge 
* No parameters

xprecharge_82 
+ vdd bl[82] br[82] en_b 
+ precharge 
* No parameters

xprecharge_83 
+ vdd bl[83] br[83] en_b 
+ precharge 
* No parameters

xprecharge_84 
+ vdd bl[84] br[84] en_b 
+ precharge 
* No parameters

xprecharge_85 
+ vdd bl[85] br[85] en_b 
+ precharge 
* No parameters

xprecharge_86 
+ vdd bl[86] br[86] en_b 
+ precharge 
* No parameters

xprecharge_87 
+ vdd bl[87] br[87] en_b 
+ precharge 
* No parameters

xprecharge_88 
+ vdd bl[88] br[88] en_b 
+ precharge 
* No parameters

xprecharge_89 
+ vdd bl[89] br[89] en_b 
+ precharge 
* No parameters

xprecharge_90 
+ vdd bl[90] br[90] en_b 
+ precharge 
* No parameters

xprecharge_91 
+ vdd bl[91] br[91] en_b 
+ precharge 
* No parameters

xprecharge_92 
+ vdd bl[92] br[92] en_b 
+ precharge 
* No parameters

xprecharge_93 
+ vdd bl[93] br[93] en_b 
+ precharge 
* No parameters

xprecharge_94 
+ vdd bl[94] br[94] en_b 
+ precharge 
* No parameters

xprecharge_95 
+ vdd bl[95] br[95] en_b 
+ precharge 
* No parameters

xprecharge_96 
+ vdd bl[96] br[96] en_b 
+ precharge 
* No parameters

xprecharge_97 
+ vdd bl[97] br[97] en_b 
+ precharge 
* No parameters

xprecharge_98 
+ vdd bl[98] br[98] en_b 
+ precharge 
* No parameters

xprecharge_99 
+ vdd bl[99] br[99] en_b 
+ precharge 
* No parameters

xprecharge_100 
+ vdd bl[100] br[100] en_b 
+ precharge 
* No parameters

xprecharge_101 
+ vdd bl[101] br[101] en_b 
+ precharge 
* No parameters

xprecharge_102 
+ vdd bl[102] br[102] en_b 
+ precharge 
* No parameters

xprecharge_103 
+ vdd bl[103] br[103] en_b 
+ precharge 
* No parameters

xprecharge_104 
+ vdd bl[104] br[104] en_b 
+ precharge 
* No parameters

xprecharge_105 
+ vdd bl[105] br[105] en_b 
+ precharge 
* No parameters

xprecharge_106 
+ vdd bl[106] br[106] en_b 
+ precharge 
* No parameters

xprecharge_107 
+ vdd bl[107] br[107] en_b 
+ precharge 
* No parameters

xprecharge_108 
+ vdd bl[108] br[108] en_b 
+ precharge 
* No parameters

xprecharge_109 
+ vdd bl[109] br[109] en_b 
+ precharge 
* No parameters

xprecharge_110 
+ vdd bl[110] br[110] en_b 
+ precharge 
* No parameters

xprecharge_111 
+ vdd bl[111] br[111] en_b 
+ precharge 
* No parameters

xprecharge_112 
+ vdd bl[112] br[112] en_b 
+ precharge 
* No parameters

xprecharge_113 
+ vdd bl[113] br[113] en_b 
+ precharge 
* No parameters

xprecharge_114 
+ vdd bl[114] br[114] en_b 
+ precharge 
* No parameters

xprecharge_115 
+ vdd bl[115] br[115] en_b 
+ precharge 
* No parameters

xprecharge_116 
+ vdd bl[116] br[116] en_b 
+ precharge 
* No parameters

xprecharge_117 
+ vdd bl[117] br[117] en_b 
+ precharge 
* No parameters

xprecharge_118 
+ vdd bl[118] br[118] en_b 
+ precharge 
* No parameters

xprecharge_119 
+ vdd bl[119] br[119] en_b 
+ precharge 
* No parameters

xprecharge_120 
+ vdd bl[120] br[120] en_b 
+ precharge 
* No parameters

xprecharge_121 
+ vdd bl[121] br[121] en_b 
+ precharge 
* No parameters

xprecharge_122 
+ vdd bl[122] br[122] en_b 
+ precharge 
* No parameters

xprecharge_123 
+ vdd bl[123] br[123] en_b 
+ precharge 
* No parameters

xprecharge_124 
+ vdd bl[124] br[124] en_b 
+ precharge 
* No parameters

xprecharge_125 
+ vdd bl[125] br[125] en_b 
+ precharge 
* No parameters

xprecharge_126 
+ vdd bl[126] br[126] en_b 
+ precharge 
* No parameters

xprecharge_127 
+ vdd bl[127] br[127] en_b 
+ precharge 
* No parameters

xprecharge_128 
+ vdd bl[128] br[128] en_b 
+ precharge 
* No parameters

.ENDS

.SUBCKT read_mux 
+ sel_b bl br bl_out br_out vdd 

xMBL 
+ bl_out sel_b bl vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

xMBR 
+ br_out sel_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

.ENDS

.SUBCKT read_mux_array 
+ sel_b[1] sel_b[0] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_out[63] bl_out[62] bl_out[61] bl_out[60] bl_out[59] bl_out[58] bl_out[57] bl_out[56] bl_out[55] bl_out[54] bl_out[53] bl_out[52] bl_out[51] bl_out[50] bl_out[49] bl_out[48] bl_out[47] bl_out[46] bl_out[45] bl_out[44] bl_out[43] bl_out[42] bl_out[41] bl_out[40] bl_out[39] bl_out[38] bl_out[37] bl_out[36] bl_out[35] bl_out[34] bl_out[33] bl_out[32] bl_out[31] bl_out[30] bl_out[29] bl_out[28] bl_out[27] bl_out[26] bl_out[25] bl_out[24] bl_out[23] bl_out[22] bl_out[21] bl_out[20] bl_out[19] bl_out[18] bl_out[17] bl_out[16] bl_out[15] bl_out[14] bl_out[13] bl_out[12] bl_out[11] bl_out[10] bl_out[9] bl_out[8] bl_out[7] bl_out[6] bl_out[5] bl_out[4] bl_out[3] bl_out[2] bl_out[1] bl_out[0] br_out[63] br_out[62] br_out[61] br_out[60] br_out[59] br_out[58] br_out[57] br_out[56] br_out[55] br_out[54] br_out[53] br_out[52] br_out[51] br_out[50] br_out[49] br_out[48] br_out[47] br_out[46] br_out[45] br_out[44] br_out[43] br_out[42] br_out[41] br_out[40] br_out[39] br_out[38] br_out[37] br_out[36] br_out[35] br_out[34] br_out[33] br_out[32] br_out[31] br_out[30] br_out[29] br_out[28] br_out[27] br_out[26] br_out[25] br_out[24] br_out[23] br_out[22] br_out[21] br_out[20] br_out[19] br_out[18] br_out[17] br_out[16] br_out[15] br_out[14] br_out[13] br_out[12] br_out[11] br_out[10] br_out[9] br_out[8] br_out[7] br_out[6] br_out[5] br_out[4] br_out[3] br_out[2] br_out[1] br_out[0] vdd 

xmux_0 
+ sel_b[0] bl[0] br[0] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_1 
+ sel_b[1] bl[1] br[1] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_2 
+ sel_b[0] bl[2] br[2] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_3 
+ sel_b[1] bl[3] br[3] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_4 
+ sel_b[0] bl[4] br[4] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_5 
+ sel_b[1] bl[5] br[5] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_6 
+ sel_b[0] bl[6] br[6] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_7 
+ sel_b[1] bl[7] br[7] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_8 
+ sel_b[0] bl[8] br[8] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_9 
+ sel_b[1] bl[9] br[9] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_10 
+ sel_b[0] bl[10] br[10] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_11 
+ sel_b[1] bl[11] br[11] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_12 
+ sel_b[0] bl[12] br[12] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_13 
+ sel_b[1] bl[13] br[13] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_14 
+ sel_b[0] bl[14] br[14] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_15 
+ sel_b[1] bl[15] br[15] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_16 
+ sel_b[0] bl[16] br[16] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_17 
+ sel_b[1] bl[17] br[17] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_18 
+ sel_b[0] bl[18] br[18] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_19 
+ sel_b[1] bl[19] br[19] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_20 
+ sel_b[0] bl[20] br[20] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_21 
+ sel_b[1] bl[21] br[21] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_22 
+ sel_b[0] bl[22] br[22] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_23 
+ sel_b[1] bl[23] br[23] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_24 
+ sel_b[0] bl[24] br[24] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_25 
+ sel_b[1] bl[25] br[25] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_26 
+ sel_b[0] bl[26] br[26] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_27 
+ sel_b[1] bl[27] br[27] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_28 
+ sel_b[0] bl[28] br[28] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_29 
+ sel_b[1] bl[29] br[29] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_30 
+ sel_b[0] bl[30] br[30] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_31 
+ sel_b[1] bl[31] br[31] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_32 
+ sel_b[0] bl[32] br[32] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_33 
+ sel_b[1] bl[33] br[33] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_34 
+ sel_b[0] bl[34] br[34] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_35 
+ sel_b[1] bl[35] br[35] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_36 
+ sel_b[0] bl[36] br[36] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_37 
+ sel_b[1] bl[37] br[37] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_38 
+ sel_b[0] bl[38] br[38] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_39 
+ sel_b[1] bl[39] br[39] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_40 
+ sel_b[0] bl[40] br[40] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_41 
+ sel_b[1] bl[41] br[41] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_42 
+ sel_b[0] bl[42] br[42] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_43 
+ sel_b[1] bl[43] br[43] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_44 
+ sel_b[0] bl[44] br[44] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_45 
+ sel_b[1] bl[45] br[45] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_46 
+ sel_b[0] bl[46] br[46] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_47 
+ sel_b[1] bl[47] br[47] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_48 
+ sel_b[0] bl[48] br[48] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_49 
+ sel_b[1] bl[49] br[49] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_50 
+ sel_b[0] bl[50] br[50] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_51 
+ sel_b[1] bl[51] br[51] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_52 
+ sel_b[0] bl[52] br[52] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_53 
+ sel_b[1] bl[53] br[53] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_54 
+ sel_b[0] bl[54] br[54] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_55 
+ sel_b[1] bl[55] br[55] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_56 
+ sel_b[0] bl[56] br[56] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_57 
+ sel_b[1] bl[57] br[57] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_58 
+ sel_b[0] bl[58] br[58] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_59 
+ sel_b[1] bl[59] br[59] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_60 
+ sel_b[0] bl[60] br[60] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_61 
+ sel_b[1] bl[61] br[61] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_62 
+ sel_b[0] bl[62] br[62] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_63 
+ sel_b[1] bl[63] br[63] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_64 
+ sel_b[0] bl[64] br[64] bl_out[32] br_out[32] vdd 
+ read_mux 
* No parameters

xmux_65 
+ sel_b[1] bl[65] br[65] bl_out[32] br_out[32] vdd 
+ read_mux 
* No parameters

xmux_66 
+ sel_b[0] bl[66] br[66] bl_out[33] br_out[33] vdd 
+ read_mux 
* No parameters

xmux_67 
+ sel_b[1] bl[67] br[67] bl_out[33] br_out[33] vdd 
+ read_mux 
* No parameters

xmux_68 
+ sel_b[0] bl[68] br[68] bl_out[34] br_out[34] vdd 
+ read_mux 
* No parameters

xmux_69 
+ sel_b[1] bl[69] br[69] bl_out[34] br_out[34] vdd 
+ read_mux 
* No parameters

xmux_70 
+ sel_b[0] bl[70] br[70] bl_out[35] br_out[35] vdd 
+ read_mux 
* No parameters

xmux_71 
+ sel_b[1] bl[71] br[71] bl_out[35] br_out[35] vdd 
+ read_mux 
* No parameters

xmux_72 
+ sel_b[0] bl[72] br[72] bl_out[36] br_out[36] vdd 
+ read_mux 
* No parameters

xmux_73 
+ sel_b[1] bl[73] br[73] bl_out[36] br_out[36] vdd 
+ read_mux 
* No parameters

xmux_74 
+ sel_b[0] bl[74] br[74] bl_out[37] br_out[37] vdd 
+ read_mux 
* No parameters

xmux_75 
+ sel_b[1] bl[75] br[75] bl_out[37] br_out[37] vdd 
+ read_mux 
* No parameters

xmux_76 
+ sel_b[0] bl[76] br[76] bl_out[38] br_out[38] vdd 
+ read_mux 
* No parameters

xmux_77 
+ sel_b[1] bl[77] br[77] bl_out[38] br_out[38] vdd 
+ read_mux 
* No parameters

xmux_78 
+ sel_b[0] bl[78] br[78] bl_out[39] br_out[39] vdd 
+ read_mux 
* No parameters

xmux_79 
+ sel_b[1] bl[79] br[79] bl_out[39] br_out[39] vdd 
+ read_mux 
* No parameters

xmux_80 
+ sel_b[0] bl[80] br[80] bl_out[40] br_out[40] vdd 
+ read_mux 
* No parameters

xmux_81 
+ sel_b[1] bl[81] br[81] bl_out[40] br_out[40] vdd 
+ read_mux 
* No parameters

xmux_82 
+ sel_b[0] bl[82] br[82] bl_out[41] br_out[41] vdd 
+ read_mux 
* No parameters

xmux_83 
+ sel_b[1] bl[83] br[83] bl_out[41] br_out[41] vdd 
+ read_mux 
* No parameters

xmux_84 
+ sel_b[0] bl[84] br[84] bl_out[42] br_out[42] vdd 
+ read_mux 
* No parameters

xmux_85 
+ sel_b[1] bl[85] br[85] bl_out[42] br_out[42] vdd 
+ read_mux 
* No parameters

xmux_86 
+ sel_b[0] bl[86] br[86] bl_out[43] br_out[43] vdd 
+ read_mux 
* No parameters

xmux_87 
+ sel_b[1] bl[87] br[87] bl_out[43] br_out[43] vdd 
+ read_mux 
* No parameters

xmux_88 
+ sel_b[0] bl[88] br[88] bl_out[44] br_out[44] vdd 
+ read_mux 
* No parameters

xmux_89 
+ sel_b[1] bl[89] br[89] bl_out[44] br_out[44] vdd 
+ read_mux 
* No parameters

xmux_90 
+ sel_b[0] bl[90] br[90] bl_out[45] br_out[45] vdd 
+ read_mux 
* No parameters

xmux_91 
+ sel_b[1] bl[91] br[91] bl_out[45] br_out[45] vdd 
+ read_mux 
* No parameters

xmux_92 
+ sel_b[0] bl[92] br[92] bl_out[46] br_out[46] vdd 
+ read_mux 
* No parameters

xmux_93 
+ sel_b[1] bl[93] br[93] bl_out[46] br_out[46] vdd 
+ read_mux 
* No parameters

xmux_94 
+ sel_b[0] bl[94] br[94] bl_out[47] br_out[47] vdd 
+ read_mux 
* No parameters

xmux_95 
+ sel_b[1] bl[95] br[95] bl_out[47] br_out[47] vdd 
+ read_mux 
* No parameters

xmux_96 
+ sel_b[0] bl[96] br[96] bl_out[48] br_out[48] vdd 
+ read_mux 
* No parameters

xmux_97 
+ sel_b[1] bl[97] br[97] bl_out[48] br_out[48] vdd 
+ read_mux 
* No parameters

xmux_98 
+ sel_b[0] bl[98] br[98] bl_out[49] br_out[49] vdd 
+ read_mux 
* No parameters

xmux_99 
+ sel_b[1] bl[99] br[99] bl_out[49] br_out[49] vdd 
+ read_mux 
* No parameters

xmux_100 
+ sel_b[0] bl[100] br[100] bl_out[50] br_out[50] vdd 
+ read_mux 
* No parameters

xmux_101 
+ sel_b[1] bl[101] br[101] bl_out[50] br_out[50] vdd 
+ read_mux 
* No parameters

xmux_102 
+ sel_b[0] bl[102] br[102] bl_out[51] br_out[51] vdd 
+ read_mux 
* No parameters

xmux_103 
+ sel_b[1] bl[103] br[103] bl_out[51] br_out[51] vdd 
+ read_mux 
* No parameters

xmux_104 
+ sel_b[0] bl[104] br[104] bl_out[52] br_out[52] vdd 
+ read_mux 
* No parameters

xmux_105 
+ sel_b[1] bl[105] br[105] bl_out[52] br_out[52] vdd 
+ read_mux 
* No parameters

xmux_106 
+ sel_b[0] bl[106] br[106] bl_out[53] br_out[53] vdd 
+ read_mux 
* No parameters

xmux_107 
+ sel_b[1] bl[107] br[107] bl_out[53] br_out[53] vdd 
+ read_mux 
* No parameters

xmux_108 
+ sel_b[0] bl[108] br[108] bl_out[54] br_out[54] vdd 
+ read_mux 
* No parameters

xmux_109 
+ sel_b[1] bl[109] br[109] bl_out[54] br_out[54] vdd 
+ read_mux 
* No parameters

xmux_110 
+ sel_b[0] bl[110] br[110] bl_out[55] br_out[55] vdd 
+ read_mux 
* No parameters

xmux_111 
+ sel_b[1] bl[111] br[111] bl_out[55] br_out[55] vdd 
+ read_mux 
* No parameters

xmux_112 
+ sel_b[0] bl[112] br[112] bl_out[56] br_out[56] vdd 
+ read_mux 
* No parameters

xmux_113 
+ sel_b[1] bl[113] br[113] bl_out[56] br_out[56] vdd 
+ read_mux 
* No parameters

xmux_114 
+ sel_b[0] bl[114] br[114] bl_out[57] br_out[57] vdd 
+ read_mux 
* No parameters

xmux_115 
+ sel_b[1] bl[115] br[115] bl_out[57] br_out[57] vdd 
+ read_mux 
* No parameters

xmux_116 
+ sel_b[0] bl[116] br[116] bl_out[58] br_out[58] vdd 
+ read_mux 
* No parameters

xmux_117 
+ sel_b[1] bl[117] br[117] bl_out[58] br_out[58] vdd 
+ read_mux 
* No parameters

xmux_118 
+ sel_b[0] bl[118] br[118] bl_out[59] br_out[59] vdd 
+ read_mux 
* No parameters

xmux_119 
+ sel_b[1] bl[119] br[119] bl_out[59] br_out[59] vdd 
+ read_mux 
* No parameters

xmux_120 
+ sel_b[0] bl[120] br[120] bl_out[60] br_out[60] vdd 
+ read_mux 
* No parameters

xmux_121 
+ sel_b[1] bl[121] br[121] bl_out[60] br_out[60] vdd 
+ read_mux 
* No parameters

xmux_122 
+ sel_b[0] bl[122] br[122] bl_out[61] br_out[61] vdd 
+ read_mux 
* No parameters

xmux_123 
+ sel_b[1] bl[123] br[123] bl_out[61] br_out[61] vdd 
+ read_mux 
* No parameters

xmux_124 
+ sel_b[0] bl[124] br[124] bl_out[62] br_out[62] vdd 
+ read_mux 
* No parameters

xmux_125 
+ sel_b[1] bl[125] br[125] bl_out[62] br_out[62] vdd 
+ read_mux 
* No parameters

xmux_126 
+ sel_b[0] bl[126] br[126] bl_out[63] br_out[63] vdd 
+ read_mux 
* No parameters

xmux_127 
+ sel_b[1] bl[127] br[127] bl_out[63] br_out[63] vdd 
+ read_mux 
* No parameters

.ENDS

.SUBCKT write_mux 
+ we data data_b bl br vss 

xMMUXBR 
+ br data x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMMUXBL 
+ bl data_b x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMPD 
+ x we vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT write_mux_array 
+ we[1] we[0] data[63] data[62] data[61] data[60] data[59] data[58] data[57] data[56] data[55] data[54] data[53] data[52] data[51] data[50] data[49] data[48] data[47] data[46] data[45] data[44] data[43] data[42] data[41] data[40] data[39] data[38] data[37] data[36] data[35] data[34] data[33] data[32] data[31] data[30] data[29] data[28] data[27] data[26] data[25] data[24] data[23] data[22] data[21] data[20] data[19] data[18] data[17] data[16] data[15] data[14] data[13] data[12] data[11] data[10] data[9] data[8] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[63] data_b[62] data_b[61] data_b[60] data_b[59] data_b[58] data_b[57] data_b[56] data_b[55] data_b[54] data_b[53] data_b[52] data_b[51] data_b[50] data_b[49] data_b[48] data_b[47] data_b[46] data_b[45] data_b[44] data_b[43] data_b[42] data_b[41] data_b[40] data_b[39] data_b[38] data_b[37] data_b[36] data_b[35] data_b[34] data_b[33] data_b[32] data_b[31] data_b[30] data_b[29] data_b[28] data_b[27] data_b[26] data_b[25] data_b[24] data_b[23] data_b[22] data_b[21] data_b[20] data_b[19] data_b[18] data_b[17] data_b[16] data_b[15] data_b[14] data_b[13] data_b[12] data_b[11] data_b[10] data_b[9] data_b[8] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 

xmux_0 
+ we[0] data[0] data_b[0] bl[0] br[0] vss 
+ write_mux 
* No parameters

xmux_1 
+ we[1] data[0] data_b[0] bl[1] br[1] vss 
+ write_mux 
* No parameters

xmux_2 
+ we[0] data[1] data_b[1] bl[2] br[2] vss 
+ write_mux 
* No parameters

xmux_3 
+ we[1] data[1] data_b[1] bl[3] br[3] vss 
+ write_mux 
* No parameters

xmux_4 
+ we[0] data[2] data_b[2] bl[4] br[4] vss 
+ write_mux 
* No parameters

xmux_5 
+ we[1] data[2] data_b[2] bl[5] br[5] vss 
+ write_mux 
* No parameters

xmux_6 
+ we[0] data[3] data_b[3] bl[6] br[6] vss 
+ write_mux 
* No parameters

xmux_7 
+ we[1] data[3] data_b[3] bl[7] br[7] vss 
+ write_mux 
* No parameters

xmux_8 
+ we[0] data[4] data_b[4] bl[8] br[8] vss 
+ write_mux 
* No parameters

xmux_9 
+ we[1] data[4] data_b[4] bl[9] br[9] vss 
+ write_mux 
* No parameters

xmux_10 
+ we[0] data[5] data_b[5] bl[10] br[10] vss 
+ write_mux 
* No parameters

xmux_11 
+ we[1] data[5] data_b[5] bl[11] br[11] vss 
+ write_mux 
* No parameters

xmux_12 
+ we[0] data[6] data_b[6] bl[12] br[12] vss 
+ write_mux 
* No parameters

xmux_13 
+ we[1] data[6] data_b[6] bl[13] br[13] vss 
+ write_mux 
* No parameters

xmux_14 
+ we[0] data[7] data_b[7] bl[14] br[14] vss 
+ write_mux 
* No parameters

xmux_15 
+ we[1] data[7] data_b[7] bl[15] br[15] vss 
+ write_mux 
* No parameters

xmux_16 
+ we[0] data[8] data_b[8] bl[16] br[16] vss 
+ write_mux 
* No parameters

xmux_17 
+ we[1] data[8] data_b[8] bl[17] br[17] vss 
+ write_mux 
* No parameters

xmux_18 
+ we[0] data[9] data_b[9] bl[18] br[18] vss 
+ write_mux 
* No parameters

xmux_19 
+ we[1] data[9] data_b[9] bl[19] br[19] vss 
+ write_mux 
* No parameters

xmux_20 
+ we[0] data[10] data_b[10] bl[20] br[20] vss 
+ write_mux 
* No parameters

xmux_21 
+ we[1] data[10] data_b[10] bl[21] br[21] vss 
+ write_mux 
* No parameters

xmux_22 
+ we[0] data[11] data_b[11] bl[22] br[22] vss 
+ write_mux 
* No parameters

xmux_23 
+ we[1] data[11] data_b[11] bl[23] br[23] vss 
+ write_mux 
* No parameters

xmux_24 
+ we[0] data[12] data_b[12] bl[24] br[24] vss 
+ write_mux 
* No parameters

xmux_25 
+ we[1] data[12] data_b[12] bl[25] br[25] vss 
+ write_mux 
* No parameters

xmux_26 
+ we[0] data[13] data_b[13] bl[26] br[26] vss 
+ write_mux 
* No parameters

xmux_27 
+ we[1] data[13] data_b[13] bl[27] br[27] vss 
+ write_mux 
* No parameters

xmux_28 
+ we[0] data[14] data_b[14] bl[28] br[28] vss 
+ write_mux 
* No parameters

xmux_29 
+ we[1] data[14] data_b[14] bl[29] br[29] vss 
+ write_mux 
* No parameters

xmux_30 
+ we[0] data[15] data_b[15] bl[30] br[30] vss 
+ write_mux 
* No parameters

xmux_31 
+ we[1] data[15] data_b[15] bl[31] br[31] vss 
+ write_mux 
* No parameters

xmux_32 
+ we[0] data[16] data_b[16] bl[32] br[32] vss 
+ write_mux 
* No parameters

xmux_33 
+ we[1] data[16] data_b[16] bl[33] br[33] vss 
+ write_mux 
* No parameters

xmux_34 
+ we[0] data[17] data_b[17] bl[34] br[34] vss 
+ write_mux 
* No parameters

xmux_35 
+ we[1] data[17] data_b[17] bl[35] br[35] vss 
+ write_mux 
* No parameters

xmux_36 
+ we[0] data[18] data_b[18] bl[36] br[36] vss 
+ write_mux 
* No parameters

xmux_37 
+ we[1] data[18] data_b[18] bl[37] br[37] vss 
+ write_mux 
* No parameters

xmux_38 
+ we[0] data[19] data_b[19] bl[38] br[38] vss 
+ write_mux 
* No parameters

xmux_39 
+ we[1] data[19] data_b[19] bl[39] br[39] vss 
+ write_mux 
* No parameters

xmux_40 
+ we[0] data[20] data_b[20] bl[40] br[40] vss 
+ write_mux 
* No parameters

xmux_41 
+ we[1] data[20] data_b[20] bl[41] br[41] vss 
+ write_mux 
* No parameters

xmux_42 
+ we[0] data[21] data_b[21] bl[42] br[42] vss 
+ write_mux 
* No parameters

xmux_43 
+ we[1] data[21] data_b[21] bl[43] br[43] vss 
+ write_mux 
* No parameters

xmux_44 
+ we[0] data[22] data_b[22] bl[44] br[44] vss 
+ write_mux 
* No parameters

xmux_45 
+ we[1] data[22] data_b[22] bl[45] br[45] vss 
+ write_mux 
* No parameters

xmux_46 
+ we[0] data[23] data_b[23] bl[46] br[46] vss 
+ write_mux 
* No parameters

xmux_47 
+ we[1] data[23] data_b[23] bl[47] br[47] vss 
+ write_mux 
* No parameters

xmux_48 
+ we[0] data[24] data_b[24] bl[48] br[48] vss 
+ write_mux 
* No parameters

xmux_49 
+ we[1] data[24] data_b[24] bl[49] br[49] vss 
+ write_mux 
* No parameters

xmux_50 
+ we[0] data[25] data_b[25] bl[50] br[50] vss 
+ write_mux 
* No parameters

xmux_51 
+ we[1] data[25] data_b[25] bl[51] br[51] vss 
+ write_mux 
* No parameters

xmux_52 
+ we[0] data[26] data_b[26] bl[52] br[52] vss 
+ write_mux 
* No parameters

xmux_53 
+ we[1] data[26] data_b[26] bl[53] br[53] vss 
+ write_mux 
* No parameters

xmux_54 
+ we[0] data[27] data_b[27] bl[54] br[54] vss 
+ write_mux 
* No parameters

xmux_55 
+ we[1] data[27] data_b[27] bl[55] br[55] vss 
+ write_mux 
* No parameters

xmux_56 
+ we[0] data[28] data_b[28] bl[56] br[56] vss 
+ write_mux 
* No parameters

xmux_57 
+ we[1] data[28] data_b[28] bl[57] br[57] vss 
+ write_mux 
* No parameters

xmux_58 
+ we[0] data[29] data_b[29] bl[58] br[58] vss 
+ write_mux 
* No parameters

xmux_59 
+ we[1] data[29] data_b[29] bl[59] br[59] vss 
+ write_mux 
* No parameters

xmux_60 
+ we[0] data[30] data_b[30] bl[60] br[60] vss 
+ write_mux 
* No parameters

xmux_61 
+ we[1] data[30] data_b[30] bl[61] br[61] vss 
+ write_mux 
* No parameters

xmux_62 
+ we[0] data[31] data_b[31] bl[62] br[62] vss 
+ write_mux 
* No parameters

xmux_63 
+ we[1] data[31] data_b[31] bl[63] br[63] vss 
+ write_mux 
* No parameters

xmux_64 
+ we[0] data[32] data_b[32] bl[64] br[64] vss 
+ write_mux 
* No parameters

xmux_65 
+ we[1] data[32] data_b[32] bl[65] br[65] vss 
+ write_mux 
* No parameters

xmux_66 
+ we[0] data[33] data_b[33] bl[66] br[66] vss 
+ write_mux 
* No parameters

xmux_67 
+ we[1] data[33] data_b[33] bl[67] br[67] vss 
+ write_mux 
* No parameters

xmux_68 
+ we[0] data[34] data_b[34] bl[68] br[68] vss 
+ write_mux 
* No parameters

xmux_69 
+ we[1] data[34] data_b[34] bl[69] br[69] vss 
+ write_mux 
* No parameters

xmux_70 
+ we[0] data[35] data_b[35] bl[70] br[70] vss 
+ write_mux 
* No parameters

xmux_71 
+ we[1] data[35] data_b[35] bl[71] br[71] vss 
+ write_mux 
* No parameters

xmux_72 
+ we[0] data[36] data_b[36] bl[72] br[72] vss 
+ write_mux 
* No parameters

xmux_73 
+ we[1] data[36] data_b[36] bl[73] br[73] vss 
+ write_mux 
* No parameters

xmux_74 
+ we[0] data[37] data_b[37] bl[74] br[74] vss 
+ write_mux 
* No parameters

xmux_75 
+ we[1] data[37] data_b[37] bl[75] br[75] vss 
+ write_mux 
* No parameters

xmux_76 
+ we[0] data[38] data_b[38] bl[76] br[76] vss 
+ write_mux 
* No parameters

xmux_77 
+ we[1] data[38] data_b[38] bl[77] br[77] vss 
+ write_mux 
* No parameters

xmux_78 
+ we[0] data[39] data_b[39] bl[78] br[78] vss 
+ write_mux 
* No parameters

xmux_79 
+ we[1] data[39] data_b[39] bl[79] br[79] vss 
+ write_mux 
* No parameters

xmux_80 
+ we[0] data[40] data_b[40] bl[80] br[80] vss 
+ write_mux 
* No parameters

xmux_81 
+ we[1] data[40] data_b[40] bl[81] br[81] vss 
+ write_mux 
* No parameters

xmux_82 
+ we[0] data[41] data_b[41] bl[82] br[82] vss 
+ write_mux 
* No parameters

xmux_83 
+ we[1] data[41] data_b[41] bl[83] br[83] vss 
+ write_mux 
* No parameters

xmux_84 
+ we[0] data[42] data_b[42] bl[84] br[84] vss 
+ write_mux 
* No parameters

xmux_85 
+ we[1] data[42] data_b[42] bl[85] br[85] vss 
+ write_mux 
* No parameters

xmux_86 
+ we[0] data[43] data_b[43] bl[86] br[86] vss 
+ write_mux 
* No parameters

xmux_87 
+ we[1] data[43] data_b[43] bl[87] br[87] vss 
+ write_mux 
* No parameters

xmux_88 
+ we[0] data[44] data_b[44] bl[88] br[88] vss 
+ write_mux 
* No parameters

xmux_89 
+ we[1] data[44] data_b[44] bl[89] br[89] vss 
+ write_mux 
* No parameters

xmux_90 
+ we[0] data[45] data_b[45] bl[90] br[90] vss 
+ write_mux 
* No parameters

xmux_91 
+ we[1] data[45] data_b[45] bl[91] br[91] vss 
+ write_mux 
* No parameters

xmux_92 
+ we[0] data[46] data_b[46] bl[92] br[92] vss 
+ write_mux 
* No parameters

xmux_93 
+ we[1] data[46] data_b[46] bl[93] br[93] vss 
+ write_mux 
* No parameters

xmux_94 
+ we[0] data[47] data_b[47] bl[94] br[94] vss 
+ write_mux 
* No parameters

xmux_95 
+ we[1] data[47] data_b[47] bl[95] br[95] vss 
+ write_mux 
* No parameters

xmux_96 
+ we[0] data[48] data_b[48] bl[96] br[96] vss 
+ write_mux 
* No parameters

xmux_97 
+ we[1] data[48] data_b[48] bl[97] br[97] vss 
+ write_mux 
* No parameters

xmux_98 
+ we[0] data[49] data_b[49] bl[98] br[98] vss 
+ write_mux 
* No parameters

xmux_99 
+ we[1] data[49] data_b[49] bl[99] br[99] vss 
+ write_mux 
* No parameters

xmux_100 
+ we[0] data[50] data_b[50] bl[100] br[100] vss 
+ write_mux 
* No parameters

xmux_101 
+ we[1] data[50] data_b[50] bl[101] br[101] vss 
+ write_mux 
* No parameters

xmux_102 
+ we[0] data[51] data_b[51] bl[102] br[102] vss 
+ write_mux 
* No parameters

xmux_103 
+ we[1] data[51] data_b[51] bl[103] br[103] vss 
+ write_mux 
* No parameters

xmux_104 
+ we[0] data[52] data_b[52] bl[104] br[104] vss 
+ write_mux 
* No parameters

xmux_105 
+ we[1] data[52] data_b[52] bl[105] br[105] vss 
+ write_mux 
* No parameters

xmux_106 
+ we[0] data[53] data_b[53] bl[106] br[106] vss 
+ write_mux 
* No parameters

xmux_107 
+ we[1] data[53] data_b[53] bl[107] br[107] vss 
+ write_mux 
* No parameters

xmux_108 
+ we[0] data[54] data_b[54] bl[108] br[108] vss 
+ write_mux 
* No parameters

xmux_109 
+ we[1] data[54] data_b[54] bl[109] br[109] vss 
+ write_mux 
* No parameters

xmux_110 
+ we[0] data[55] data_b[55] bl[110] br[110] vss 
+ write_mux 
* No parameters

xmux_111 
+ we[1] data[55] data_b[55] bl[111] br[111] vss 
+ write_mux 
* No parameters

xmux_112 
+ we[0] data[56] data_b[56] bl[112] br[112] vss 
+ write_mux 
* No parameters

xmux_113 
+ we[1] data[56] data_b[56] bl[113] br[113] vss 
+ write_mux 
* No parameters

xmux_114 
+ we[0] data[57] data_b[57] bl[114] br[114] vss 
+ write_mux 
* No parameters

xmux_115 
+ we[1] data[57] data_b[57] bl[115] br[115] vss 
+ write_mux 
* No parameters

xmux_116 
+ we[0] data[58] data_b[58] bl[116] br[116] vss 
+ write_mux 
* No parameters

xmux_117 
+ we[1] data[58] data_b[58] bl[117] br[117] vss 
+ write_mux 
* No parameters

xmux_118 
+ we[0] data[59] data_b[59] bl[118] br[118] vss 
+ write_mux 
* No parameters

xmux_119 
+ we[1] data[59] data_b[59] bl[119] br[119] vss 
+ write_mux 
* No parameters

xmux_120 
+ we[0] data[60] data_b[60] bl[120] br[120] vss 
+ write_mux 
* No parameters

xmux_121 
+ we[1] data[60] data_b[60] bl[121] br[121] vss 
+ write_mux 
* No parameters

xmux_122 
+ we[0] data[61] data_b[61] bl[122] br[122] vss 
+ write_mux 
* No parameters

xmux_123 
+ we[1] data[61] data_b[61] bl[123] br[123] vss 
+ write_mux 
* No parameters

xmux_124 
+ we[0] data[62] data_b[62] bl[124] br[124] vss 
+ write_mux 
* No parameters

xmux_125 
+ we[1] data[62] data_b[62] bl[125] br[125] vss 
+ write_mux 
* No parameters

xmux_126 
+ we[0] data[63] data_b[63] bl[126] br[126] vss 
+ write_mux 
* No parameters

xmux_127 
+ we[1] data[63] data_b[63] bl[127] br[127] vss 
+ write_mux 
* No parameters

.ENDS

.SUBCKT data_dff_array 
+ vdd vss clk d[63] d[62] d[61] d[60] d[59] d[58] d[57] d[56] d[55] d[54] d[53] d[52] d[51] d[50] d[49] d[48] d[47] d[46] d[45] d[44] d[43] d[42] d[41] d[40] d[39] d[38] d[37] d[36] d[35] d[34] d[33] d[32] d[31] d[30] d[29] d[28] d[27] d[26] d[25] d[24] d[23] d[22] d[21] d[20] d[19] d[18] d[17] d[16] d[15] d[14] d[13] d[12] d[11] d[10] d[9] d[8] d[7] d[6] d[5] d[4] d[3] d[2] d[1] d[0] q[63] q[62] q[61] q[60] q[59] q[58] q[57] q[56] q[55] q[54] q[53] q[52] q[51] q[50] q[49] q[48] q[47] q[46] q[45] q[44] q[43] q[42] q[41] q[40] q[39] q[38] q[37] q[36] q[35] q[34] q[33] q[32] q[31] q[30] q[29] q[28] q[27] q[26] q[25] q[24] q[23] q[22] q[21] q[20] q[19] q[18] q[17] q[16] q[15] q[14] q[13] q[12] q[11] q[10] q[9] q[8] q[7] q[6] q[5] q[4] q[3] q[2] q[1] q[0] q_b[63] q_b[62] q_b[61] q_b[60] q_b[59] q_b[58] q_b[57] q_b[56] q_b[55] q_b[54] q_b[53] q_b[52] q_b[51] q_b[50] q_b[49] q_b[48] q_b[47] q_b[46] q_b[45] q_b[44] q_b[43] q_b[42] q_b[41] q_b[40] q_b[39] q_b[38] q_b[37] q_b[36] q_b[35] q_b[34] q_b[33] q_b[32] q_b[31] q_b[30] q_b[29] q_b[28] q_b[27] q_b[26] q_b[25] q_b[24] q_b[23] q_b[22] q_b[21] q_b[20] q_b[19] q_b[18] q_b[17] q_b[16] q_b[15] q_b[14] q_b[13] q_b[12] q_b[11] q_b[10] q_b[9] q_b[8] q_b[7] q_b[6] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

xdff_6 
+ vdd vss clk d[6] q[6] q_b[6] 
+ openram_dff 
* No parameters

xdff_7 
+ vdd vss clk d[7] q[7] q_b[7] 
+ openram_dff 
* No parameters

xdff_8 
+ vdd vss clk d[8] q[8] q_b[8] 
+ openram_dff 
* No parameters

xdff_9 
+ vdd vss clk d[9] q[9] q_b[9] 
+ openram_dff 
* No parameters

xdff_10 
+ vdd vss clk d[10] q[10] q_b[10] 
+ openram_dff 
* No parameters

xdff_11 
+ vdd vss clk d[11] q[11] q_b[11] 
+ openram_dff 
* No parameters

xdff_12 
+ vdd vss clk d[12] q[12] q_b[12] 
+ openram_dff 
* No parameters

xdff_13 
+ vdd vss clk d[13] q[13] q_b[13] 
+ openram_dff 
* No parameters

xdff_14 
+ vdd vss clk d[14] q[14] q_b[14] 
+ openram_dff 
* No parameters

xdff_15 
+ vdd vss clk d[15] q[15] q_b[15] 
+ openram_dff 
* No parameters

xdff_16 
+ vdd vss clk d[16] q[16] q_b[16] 
+ openram_dff 
* No parameters

xdff_17 
+ vdd vss clk d[17] q[17] q_b[17] 
+ openram_dff 
* No parameters

xdff_18 
+ vdd vss clk d[18] q[18] q_b[18] 
+ openram_dff 
* No parameters

xdff_19 
+ vdd vss clk d[19] q[19] q_b[19] 
+ openram_dff 
* No parameters

xdff_20 
+ vdd vss clk d[20] q[20] q_b[20] 
+ openram_dff 
* No parameters

xdff_21 
+ vdd vss clk d[21] q[21] q_b[21] 
+ openram_dff 
* No parameters

xdff_22 
+ vdd vss clk d[22] q[22] q_b[22] 
+ openram_dff 
* No parameters

xdff_23 
+ vdd vss clk d[23] q[23] q_b[23] 
+ openram_dff 
* No parameters

xdff_24 
+ vdd vss clk d[24] q[24] q_b[24] 
+ openram_dff 
* No parameters

xdff_25 
+ vdd vss clk d[25] q[25] q_b[25] 
+ openram_dff 
* No parameters

xdff_26 
+ vdd vss clk d[26] q[26] q_b[26] 
+ openram_dff 
* No parameters

xdff_27 
+ vdd vss clk d[27] q[27] q_b[27] 
+ openram_dff 
* No parameters

xdff_28 
+ vdd vss clk d[28] q[28] q_b[28] 
+ openram_dff 
* No parameters

xdff_29 
+ vdd vss clk d[29] q[29] q_b[29] 
+ openram_dff 
* No parameters

xdff_30 
+ vdd vss clk d[30] q[30] q_b[30] 
+ openram_dff 
* No parameters

xdff_31 
+ vdd vss clk d[31] q[31] q_b[31] 
+ openram_dff 
* No parameters

xdff_32 
+ vdd vss clk d[32] q[32] q_b[32] 
+ openram_dff 
* No parameters

xdff_33 
+ vdd vss clk d[33] q[33] q_b[33] 
+ openram_dff 
* No parameters

xdff_34 
+ vdd vss clk d[34] q[34] q_b[34] 
+ openram_dff 
* No parameters

xdff_35 
+ vdd vss clk d[35] q[35] q_b[35] 
+ openram_dff 
* No parameters

xdff_36 
+ vdd vss clk d[36] q[36] q_b[36] 
+ openram_dff 
* No parameters

xdff_37 
+ vdd vss clk d[37] q[37] q_b[37] 
+ openram_dff 
* No parameters

xdff_38 
+ vdd vss clk d[38] q[38] q_b[38] 
+ openram_dff 
* No parameters

xdff_39 
+ vdd vss clk d[39] q[39] q_b[39] 
+ openram_dff 
* No parameters

xdff_40 
+ vdd vss clk d[40] q[40] q_b[40] 
+ openram_dff 
* No parameters

xdff_41 
+ vdd vss clk d[41] q[41] q_b[41] 
+ openram_dff 
* No parameters

xdff_42 
+ vdd vss clk d[42] q[42] q_b[42] 
+ openram_dff 
* No parameters

xdff_43 
+ vdd vss clk d[43] q[43] q_b[43] 
+ openram_dff 
* No parameters

xdff_44 
+ vdd vss clk d[44] q[44] q_b[44] 
+ openram_dff 
* No parameters

xdff_45 
+ vdd vss clk d[45] q[45] q_b[45] 
+ openram_dff 
* No parameters

xdff_46 
+ vdd vss clk d[46] q[46] q_b[46] 
+ openram_dff 
* No parameters

xdff_47 
+ vdd vss clk d[47] q[47] q_b[47] 
+ openram_dff 
* No parameters

xdff_48 
+ vdd vss clk d[48] q[48] q_b[48] 
+ openram_dff 
* No parameters

xdff_49 
+ vdd vss clk d[49] q[49] q_b[49] 
+ openram_dff 
* No parameters

xdff_50 
+ vdd vss clk d[50] q[50] q_b[50] 
+ openram_dff 
* No parameters

xdff_51 
+ vdd vss clk d[51] q[51] q_b[51] 
+ openram_dff 
* No parameters

xdff_52 
+ vdd vss clk d[52] q[52] q_b[52] 
+ openram_dff 
* No parameters

xdff_53 
+ vdd vss clk d[53] q[53] q_b[53] 
+ openram_dff 
* No parameters

xdff_54 
+ vdd vss clk d[54] q[54] q_b[54] 
+ openram_dff 
* No parameters

xdff_55 
+ vdd vss clk d[55] q[55] q_b[55] 
+ openram_dff 
* No parameters

xdff_56 
+ vdd vss clk d[56] q[56] q_b[56] 
+ openram_dff 
* No parameters

xdff_57 
+ vdd vss clk d[57] q[57] q_b[57] 
+ openram_dff 
* No parameters

xdff_58 
+ vdd vss clk d[58] q[58] q_b[58] 
+ openram_dff 
* No parameters

xdff_59 
+ vdd vss clk d[59] q[59] q_b[59] 
+ openram_dff 
* No parameters

xdff_60 
+ vdd vss clk d[60] q[60] q_b[60] 
+ openram_dff 
* No parameters

xdff_61 
+ vdd vss clk d[61] q[61] q_b[61] 
+ openram_dff 
* No parameters

xdff_62 
+ vdd vss clk d[62] q[62] q_b[62] 
+ openram_dff 
* No parameters

xdff_63 
+ vdd vss clk d[63] q[63] q_b[63] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT addr_dff_array 
+ vdd vss clk d[6] d[5] d[4] d[3] d[2] d[1] d[0] q[6] q[5] q[4] q[3] q[2] q[1] q[0] q_b[6] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

xdff_6 
+ vdd vss clk d[6] q[6] q_b[6] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT col_data_inv 
+ din din_b vdd vss 

xMP0 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.6' l='0.15' 

xMN0 
+ din_b din vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.4' l='0.15' 

.ENDS

.SUBCKT col_inv_array 
+ din[63] din[62] din[61] din[60] din[59] din[58] din[57] din[56] din[55] din[54] din[53] din[52] din[51] din[50] din[49] din[48] din[47] din[46] din[45] din[44] din[43] din[42] din[41] din[40] din[39] din[38] din[37] din[36] din[35] din[34] din[33] din[32] din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] din_b[63] din_b[62] din_b[61] din_b[60] din_b[59] din_b[58] din_b[57] din_b[56] din_b[55] din_b[54] din_b[53] din_b[52] din_b[51] din_b[50] din_b[49] din_b[48] din_b[47] din_b[46] din_b[45] din_b[44] din_b[43] din_b[42] din_b[41] din_b[40] din_b[39] din_b[38] din_b[37] din_b[36] din_b[35] din_b[34] din_b[33] din_b[32] din_b[31] din_b[30] din_b[29] din_b[28] din_b[27] din_b[26] din_b[25] din_b[24] din_b[23] din_b[22] din_b[21] din_b[20] din_b[19] din_b[18] din_b[17] din_b[16] din_b[15] din_b[14] din_b[13] din_b[12] din_b[11] din_b[10] din_b[9] din_b[8] din_b[7] din_b[6] din_b[5] din_b[4] din_b[3] din_b[2] din_b[1] din_b[0] vdd vss 

xinv_0 
+ din[0] din_b[0] vdd vss 
+ col_data_inv 
* No parameters

xinv_1 
+ din[1] din_b[1] vdd vss 
+ col_data_inv 
* No parameters

xinv_2 
+ din[2] din_b[2] vdd vss 
+ col_data_inv 
* No parameters

xinv_3 
+ din[3] din_b[3] vdd vss 
+ col_data_inv 
* No parameters

xinv_4 
+ din[4] din_b[4] vdd vss 
+ col_data_inv 
* No parameters

xinv_5 
+ din[5] din_b[5] vdd vss 
+ col_data_inv 
* No parameters

xinv_6 
+ din[6] din_b[6] vdd vss 
+ col_data_inv 
* No parameters

xinv_7 
+ din[7] din_b[7] vdd vss 
+ col_data_inv 
* No parameters

xinv_8 
+ din[8] din_b[8] vdd vss 
+ col_data_inv 
* No parameters

xinv_9 
+ din[9] din_b[9] vdd vss 
+ col_data_inv 
* No parameters

xinv_10 
+ din[10] din_b[10] vdd vss 
+ col_data_inv 
* No parameters

xinv_11 
+ din[11] din_b[11] vdd vss 
+ col_data_inv 
* No parameters

xinv_12 
+ din[12] din_b[12] vdd vss 
+ col_data_inv 
* No parameters

xinv_13 
+ din[13] din_b[13] vdd vss 
+ col_data_inv 
* No parameters

xinv_14 
+ din[14] din_b[14] vdd vss 
+ col_data_inv 
* No parameters

xinv_15 
+ din[15] din_b[15] vdd vss 
+ col_data_inv 
* No parameters

xinv_16 
+ din[16] din_b[16] vdd vss 
+ col_data_inv 
* No parameters

xinv_17 
+ din[17] din_b[17] vdd vss 
+ col_data_inv 
* No parameters

xinv_18 
+ din[18] din_b[18] vdd vss 
+ col_data_inv 
* No parameters

xinv_19 
+ din[19] din_b[19] vdd vss 
+ col_data_inv 
* No parameters

xinv_20 
+ din[20] din_b[20] vdd vss 
+ col_data_inv 
* No parameters

xinv_21 
+ din[21] din_b[21] vdd vss 
+ col_data_inv 
* No parameters

xinv_22 
+ din[22] din_b[22] vdd vss 
+ col_data_inv 
* No parameters

xinv_23 
+ din[23] din_b[23] vdd vss 
+ col_data_inv 
* No parameters

xinv_24 
+ din[24] din_b[24] vdd vss 
+ col_data_inv 
* No parameters

xinv_25 
+ din[25] din_b[25] vdd vss 
+ col_data_inv 
* No parameters

xinv_26 
+ din[26] din_b[26] vdd vss 
+ col_data_inv 
* No parameters

xinv_27 
+ din[27] din_b[27] vdd vss 
+ col_data_inv 
* No parameters

xinv_28 
+ din[28] din_b[28] vdd vss 
+ col_data_inv 
* No parameters

xinv_29 
+ din[29] din_b[29] vdd vss 
+ col_data_inv 
* No parameters

xinv_30 
+ din[30] din_b[30] vdd vss 
+ col_data_inv 
* No parameters

xinv_31 
+ din[31] din_b[31] vdd vss 
+ col_data_inv 
* No parameters

xinv_32 
+ din[32] din_b[32] vdd vss 
+ col_data_inv 
* No parameters

xinv_33 
+ din[33] din_b[33] vdd vss 
+ col_data_inv 
* No parameters

xinv_34 
+ din[34] din_b[34] vdd vss 
+ col_data_inv 
* No parameters

xinv_35 
+ din[35] din_b[35] vdd vss 
+ col_data_inv 
* No parameters

xinv_36 
+ din[36] din_b[36] vdd vss 
+ col_data_inv 
* No parameters

xinv_37 
+ din[37] din_b[37] vdd vss 
+ col_data_inv 
* No parameters

xinv_38 
+ din[38] din_b[38] vdd vss 
+ col_data_inv 
* No parameters

xinv_39 
+ din[39] din_b[39] vdd vss 
+ col_data_inv 
* No parameters

xinv_40 
+ din[40] din_b[40] vdd vss 
+ col_data_inv 
* No parameters

xinv_41 
+ din[41] din_b[41] vdd vss 
+ col_data_inv 
* No parameters

xinv_42 
+ din[42] din_b[42] vdd vss 
+ col_data_inv 
* No parameters

xinv_43 
+ din[43] din_b[43] vdd vss 
+ col_data_inv 
* No parameters

xinv_44 
+ din[44] din_b[44] vdd vss 
+ col_data_inv 
* No parameters

xinv_45 
+ din[45] din_b[45] vdd vss 
+ col_data_inv 
* No parameters

xinv_46 
+ din[46] din_b[46] vdd vss 
+ col_data_inv 
* No parameters

xinv_47 
+ din[47] din_b[47] vdd vss 
+ col_data_inv 
* No parameters

xinv_48 
+ din[48] din_b[48] vdd vss 
+ col_data_inv 
* No parameters

xinv_49 
+ din[49] din_b[49] vdd vss 
+ col_data_inv 
* No parameters

xinv_50 
+ din[50] din_b[50] vdd vss 
+ col_data_inv 
* No parameters

xinv_51 
+ din[51] din_b[51] vdd vss 
+ col_data_inv 
* No parameters

xinv_52 
+ din[52] din_b[52] vdd vss 
+ col_data_inv 
* No parameters

xinv_53 
+ din[53] din_b[53] vdd vss 
+ col_data_inv 
* No parameters

xinv_54 
+ din[54] din_b[54] vdd vss 
+ col_data_inv 
* No parameters

xinv_55 
+ din[55] din_b[55] vdd vss 
+ col_data_inv 
* No parameters

xinv_56 
+ din[56] din_b[56] vdd vss 
+ col_data_inv 
* No parameters

xinv_57 
+ din[57] din_b[57] vdd vss 
+ col_data_inv 
* No parameters

xinv_58 
+ din[58] din_b[58] vdd vss 
+ col_data_inv 
* No parameters

xinv_59 
+ din[59] din_b[59] vdd vss 
+ col_data_inv 
* No parameters

xinv_60 
+ din[60] din_b[60] vdd vss 
+ col_data_inv 
* No parameters

xinv_61 
+ din[61] din_b[61] vdd vss 
+ col_data_inv 
* No parameters

xinv_62 
+ din[62] din_b[62] vdd vss 
+ col_data_inv 
* No parameters

xinv_63 
+ din[63] din_b[63] vdd vss 
+ col_data_inv 
* No parameters

.ENDS

.SUBCKT sense_amp_array 
+ vdd vss clk bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] data[63] data[62] data[61] data[60] data[59] data[58] data[57] data[56] data[55] data[54] data[53] data[52] data[51] data[50] data[49] data[48] data[47] data[46] data[45] data[44] data[43] data[42] data[41] data[40] data[39] data[38] data[37] data[36] data[35] data[34] data[33] data[32] data[31] data[30] data[29] data[28] data[27] data[26] data[25] data[24] data[23] data[22] data[21] data[20] data[19] data[18] data[17] data[16] data[15] data[14] data[13] data[12] data[11] data[10] data[9] data[8] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[63] data_b[62] data_b[61] data_b[60] data_b[59] data_b[58] data_b[57] data_b[56] data_b[55] data_b[54] data_b[53] data_b[52] data_b[51] data_b[50] data_b[49] data_b[48] data_b[47] data_b[46] data_b[45] data_b[44] data_b[43] data_b[42] data_b[41] data_b[40] data_b[39] data_b[38] data_b[37] data_b[36] data_b[35] data_b[34] data_b[33] data_b[32] data_b[31] data_b[30] data_b[29] data_b[28] data_b[27] data_b[26] data_b[25] data_b[24] data_b[23] data_b[22] data_b[21] data_b[20] data_b[19] data_b[18] data_b[17] data_b[16] data_b[15] data_b[14] data_b[13] data_b[12] data_b[11] data_b[10] data_b[9] data_b[8] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] 

xsense_amp_0 
+ clk br[0] bl[0] data_b[0] data[0] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_1 
+ clk br[1] bl[1] data_b[1] data[1] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_2 
+ clk br[2] bl[2] data_b[2] data[2] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_3 
+ clk br[3] bl[3] data_b[3] data[3] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_4 
+ clk br[4] bl[4] data_b[4] data[4] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_5 
+ clk br[5] bl[5] data_b[5] data[5] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_6 
+ clk br[6] bl[6] data_b[6] data[6] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_7 
+ clk br[7] bl[7] data_b[7] data[7] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_8 
+ clk br[8] bl[8] data_b[8] data[8] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_9 
+ clk br[9] bl[9] data_b[9] data[9] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_10 
+ clk br[10] bl[10] data_b[10] data[10] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_11 
+ clk br[11] bl[11] data_b[11] data[11] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_12 
+ clk br[12] bl[12] data_b[12] data[12] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_13 
+ clk br[13] bl[13] data_b[13] data[13] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_14 
+ clk br[14] bl[14] data_b[14] data[14] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_15 
+ clk br[15] bl[15] data_b[15] data[15] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_16 
+ clk br[16] bl[16] data_b[16] data[16] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_17 
+ clk br[17] bl[17] data_b[17] data[17] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_18 
+ clk br[18] bl[18] data_b[18] data[18] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_19 
+ clk br[19] bl[19] data_b[19] data[19] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_20 
+ clk br[20] bl[20] data_b[20] data[20] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_21 
+ clk br[21] bl[21] data_b[21] data[21] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_22 
+ clk br[22] bl[22] data_b[22] data[22] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_23 
+ clk br[23] bl[23] data_b[23] data[23] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_24 
+ clk br[24] bl[24] data_b[24] data[24] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_25 
+ clk br[25] bl[25] data_b[25] data[25] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_26 
+ clk br[26] bl[26] data_b[26] data[26] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_27 
+ clk br[27] bl[27] data_b[27] data[27] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_28 
+ clk br[28] bl[28] data_b[28] data[28] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_29 
+ clk br[29] bl[29] data_b[29] data[29] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_30 
+ clk br[30] bl[30] data_b[30] data[30] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_31 
+ clk br[31] bl[31] data_b[31] data[31] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_32 
+ clk br[32] bl[32] data_b[32] data[32] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_33 
+ clk br[33] bl[33] data_b[33] data[33] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_34 
+ clk br[34] bl[34] data_b[34] data[34] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_35 
+ clk br[35] bl[35] data_b[35] data[35] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_36 
+ clk br[36] bl[36] data_b[36] data[36] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_37 
+ clk br[37] bl[37] data_b[37] data[37] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_38 
+ clk br[38] bl[38] data_b[38] data[38] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_39 
+ clk br[39] bl[39] data_b[39] data[39] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_40 
+ clk br[40] bl[40] data_b[40] data[40] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_41 
+ clk br[41] bl[41] data_b[41] data[41] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_42 
+ clk br[42] bl[42] data_b[42] data[42] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_43 
+ clk br[43] bl[43] data_b[43] data[43] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_44 
+ clk br[44] bl[44] data_b[44] data[44] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_45 
+ clk br[45] bl[45] data_b[45] data[45] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_46 
+ clk br[46] bl[46] data_b[46] data[46] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_47 
+ clk br[47] bl[47] data_b[47] data[47] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_48 
+ clk br[48] bl[48] data_b[48] data[48] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_49 
+ clk br[49] bl[49] data_b[49] data[49] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_50 
+ clk br[50] bl[50] data_b[50] data[50] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_51 
+ clk br[51] bl[51] data_b[51] data[51] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_52 
+ clk br[52] bl[52] data_b[52] data[52] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_53 
+ clk br[53] bl[53] data_b[53] data[53] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_54 
+ clk br[54] bl[54] data_b[54] data[54] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_55 
+ clk br[55] bl[55] data_b[55] data[55] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_56 
+ clk br[56] bl[56] data_b[56] data[56] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_57 
+ clk br[57] bl[57] data_b[57] data[57] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_58 
+ clk br[58] bl[58] data_b[58] data[58] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_59 
+ clk br[59] bl[59] data_b[59] data[59] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_60 
+ clk br[60] bl[60] data_b[60] data[60] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_61 
+ clk br[61] bl[61] data_b[61] data[61] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_62 
+ clk br[62] bl[62] data_b[62] data[62] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_63 
+ clk br[63] bl[63] data_b[63] data[63] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

.ENDS

.SUBCKT dout_buf 
+ din1 din2 dout1 dout2 vdd vss 

xMP11 
+ x1 din1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN11 
+ x1 din1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP21 
+ dout1 x1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN21 
+ dout1 x1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMP12 
+ x2 din2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN12 
+ x2 din2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP22 
+ dout2 x2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN22 
+ dout2 x2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT dout_buf_array 
+ din1[63] din1[62] din1[61] din1[60] din1[59] din1[58] din1[57] din1[56] din1[55] din1[54] din1[53] din1[52] din1[51] din1[50] din1[49] din1[48] din1[47] din1[46] din1[45] din1[44] din1[43] din1[42] din1[41] din1[40] din1[39] din1[38] din1[37] din1[36] din1[35] din1[34] din1[33] din1[32] din1[31] din1[30] din1[29] din1[28] din1[27] din1[26] din1[25] din1[24] din1[23] din1[22] din1[21] din1[20] din1[19] din1[18] din1[17] din1[16] din1[15] din1[14] din1[13] din1[12] din1[11] din1[10] din1[9] din1[8] din1[7] din1[6] din1[5] din1[4] din1[3] din1[2] din1[1] din1[0] din2[63] din2[62] din2[61] din2[60] din2[59] din2[58] din2[57] din2[56] din2[55] din2[54] din2[53] din2[52] din2[51] din2[50] din2[49] din2[48] din2[47] din2[46] din2[45] din2[44] din2[43] din2[42] din2[41] din2[40] din2[39] din2[38] din2[37] din2[36] din2[35] din2[34] din2[33] din2[32] din2[31] din2[30] din2[29] din2[28] din2[27] din2[26] din2[25] din2[24] din2[23] din2[22] din2[21] din2[20] din2[19] din2[18] din2[17] din2[16] din2[15] din2[14] din2[13] din2[12] din2[11] din2[10] din2[9] din2[8] din2[7] din2[6] din2[5] din2[4] din2[3] din2[2] din2[1] din2[0] dout1[63] dout1[62] dout1[61] dout1[60] dout1[59] dout1[58] dout1[57] dout1[56] dout1[55] dout1[54] dout1[53] dout1[52] dout1[51] dout1[50] dout1[49] dout1[48] dout1[47] dout1[46] dout1[45] dout1[44] dout1[43] dout1[42] dout1[41] dout1[40] dout1[39] dout1[38] dout1[37] dout1[36] dout1[35] dout1[34] dout1[33] dout1[32] dout1[31] dout1[30] dout1[29] dout1[28] dout1[27] dout1[26] dout1[25] dout1[24] dout1[23] dout1[22] dout1[21] dout1[20] dout1[19] dout1[18] dout1[17] dout1[16] dout1[15] dout1[14] dout1[13] dout1[12] dout1[11] dout1[10] dout1[9] dout1[8] dout1[7] dout1[6] dout1[5] dout1[4] dout1[3] dout1[2] dout1[1] dout1[0] dout2[63] dout2[62] dout2[61] dout2[60] dout2[59] dout2[58] dout2[57] dout2[56] dout2[55] dout2[54] dout2[53] dout2[52] dout2[51] dout2[50] dout2[49] dout2[48] dout2[47] dout2[46] dout2[45] dout2[44] dout2[43] dout2[42] dout2[41] dout2[40] dout2[39] dout2[38] dout2[37] dout2[36] dout2[35] dout2[34] dout2[33] dout2[32] dout2[31] dout2[30] dout2[29] dout2[28] dout2[27] dout2[26] dout2[25] dout2[24] dout2[23] dout2[22] dout2[21] dout2[20] dout2[19] dout2[18] dout2[17] dout2[16] dout2[15] dout2[14] dout2[13] dout2[12] dout2[11] dout2[10] dout2[9] dout2[8] dout2[7] dout2[6] dout2[5] dout2[4] dout2[3] dout2[2] dout2[1] dout2[0] vdd vss 

xbuf_0 
+ din1[0] din2[0] dout1[0] dout2[0] vdd vss 
+ dout_buf 
* No parameters

xbuf_1 
+ din1[1] din2[1] dout1[1] dout2[1] vdd vss 
+ dout_buf 
* No parameters

xbuf_2 
+ din1[2] din2[2] dout1[2] dout2[2] vdd vss 
+ dout_buf 
* No parameters

xbuf_3 
+ din1[3] din2[3] dout1[3] dout2[3] vdd vss 
+ dout_buf 
* No parameters

xbuf_4 
+ din1[4] din2[4] dout1[4] dout2[4] vdd vss 
+ dout_buf 
* No parameters

xbuf_5 
+ din1[5] din2[5] dout1[5] dout2[5] vdd vss 
+ dout_buf 
* No parameters

xbuf_6 
+ din1[6] din2[6] dout1[6] dout2[6] vdd vss 
+ dout_buf 
* No parameters

xbuf_7 
+ din1[7] din2[7] dout1[7] dout2[7] vdd vss 
+ dout_buf 
* No parameters

xbuf_8 
+ din1[8] din2[8] dout1[8] dout2[8] vdd vss 
+ dout_buf 
* No parameters

xbuf_9 
+ din1[9] din2[9] dout1[9] dout2[9] vdd vss 
+ dout_buf 
* No parameters

xbuf_10 
+ din1[10] din2[10] dout1[10] dout2[10] vdd vss 
+ dout_buf 
* No parameters

xbuf_11 
+ din1[11] din2[11] dout1[11] dout2[11] vdd vss 
+ dout_buf 
* No parameters

xbuf_12 
+ din1[12] din2[12] dout1[12] dout2[12] vdd vss 
+ dout_buf 
* No parameters

xbuf_13 
+ din1[13] din2[13] dout1[13] dout2[13] vdd vss 
+ dout_buf 
* No parameters

xbuf_14 
+ din1[14] din2[14] dout1[14] dout2[14] vdd vss 
+ dout_buf 
* No parameters

xbuf_15 
+ din1[15] din2[15] dout1[15] dout2[15] vdd vss 
+ dout_buf 
* No parameters

xbuf_16 
+ din1[16] din2[16] dout1[16] dout2[16] vdd vss 
+ dout_buf 
* No parameters

xbuf_17 
+ din1[17] din2[17] dout1[17] dout2[17] vdd vss 
+ dout_buf 
* No parameters

xbuf_18 
+ din1[18] din2[18] dout1[18] dout2[18] vdd vss 
+ dout_buf 
* No parameters

xbuf_19 
+ din1[19] din2[19] dout1[19] dout2[19] vdd vss 
+ dout_buf 
* No parameters

xbuf_20 
+ din1[20] din2[20] dout1[20] dout2[20] vdd vss 
+ dout_buf 
* No parameters

xbuf_21 
+ din1[21] din2[21] dout1[21] dout2[21] vdd vss 
+ dout_buf 
* No parameters

xbuf_22 
+ din1[22] din2[22] dout1[22] dout2[22] vdd vss 
+ dout_buf 
* No parameters

xbuf_23 
+ din1[23] din2[23] dout1[23] dout2[23] vdd vss 
+ dout_buf 
* No parameters

xbuf_24 
+ din1[24] din2[24] dout1[24] dout2[24] vdd vss 
+ dout_buf 
* No parameters

xbuf_25 
+ din1[25] din2[25] dout1[25] dout2[25] vdd vss 
+ dout_buf 
* No parameters

xbuf_26 
+ din1[26] din2[26] dout1[26] dout2[26] vdd vss 
+ dout_buf 
* No parameters

xbuf_27 
+ din1[27] din2[27] dout1[27] dout2[27] vdd vss 
+ dout_buf 
* No parameters

xbuf_28 
+ din1[28] din2[28] dout1[28] dout2[28] vdd vss 
+ dout_buf 
* No parameters

xbuf_29 
+ din1[29] din2[29] dout1[29] dout2[29] vdd vss 
+ dout_buf 
* No parameters

xbuf_30 
+ din1[30] din2[30] dout1[30] dout2[30] vdd vss 
+ dout_buf 
* No parameters

xbuf_31 
+ din1[31] din2[31] dout1[31] dout2[31] vdd vss 
+ dout_buf 
* No parameters

xbuf_32 
+ din1[32] din2[32] dout1[32] dout2[32] vdd vss 
+ dout_buf 
* No parameters

xbuf_33 
+ din1[33] din2[33] dout1[33] dout2[33] vdd vss 
+ dout_buf 
* No parameters

xbuf_34 
+ din1[34] din2[34] dout1[34] dout2[34] vdd vss 
+ dout_buf 
* No parameters

xbuf_35 
+ din1[35] din2[35] dout1[35] dout2[35] vdd vss 
+ dout_buf 
* No parameters

xbuf_36 
+ din1[36] din2[36] dout1[36] dout2[36] vdd vss 
+ dout_buf 
* No parameters

xbuf_37 
+ din1[37] din2[37] dout1[37] dout2[37] vdd vss 
+ dout_buf 
* No parameters

xbuf_38 
+ din1[38] din2[38] dout1[38] dout2[38] vdd vss 
+ dout_buf 
* No parameters

xbuf_39 
+ din1[39] din2[39] dout1[39] dout2[39] vdd vss 
+ dout_buf 
* No parameters

xbuf_40 
+ din1[40] din2[40] dout1[40] dout2[40] vdd vss 
+ dout_buf 
* No parameters

xbuf_41 
+ din1[41] din2[41] dout1[41] dout2[41] vdd vss 
+ dout_buf 
* No parameters

xbuf_42 
+ din1[42] din2[42] dout1[42] dout2[42] vdd vss 
+ dout_buf 
* No parameters

xbuf_43 
+ din1[43] din2[43] dout1[43] dout2[43] vdd vss 
+ dout_buf 
* No parameters

xbuf_44 
+ din1[44] din2[44] dout1[44] dout2[44] vdd vss 
+ dout_buf 
* No parameters

xbuf_45 
+ din1[45] din2[45] dout1[45] dout2[45] vdd vss 
+ dout_buf 
* No parameters

xbuf_46 
+ din1[46] din2[46] dout1[46] dout2[46] vdd vss 
+ dout_buf 
* No parameters

xbuf_47 
+ din1[47] din2[47] dout1[47] dout2[47] vdd vss 
+ dout_buf 
* No parameters

xbuf_48 
+ din1[48] din2[48] dout1[48] dout2[48] vdd vss 
+ dout_buf 
* No parameters

xbuf_49 
+ din1[49] din2[49] dout1[49] dout2[49] vdd vss 
+ dout_buf 
* No parameters

xbuf_50 
+ din1[50] din2[50] dout1[50] dout2[50] vdd vss 
+ dout_buf 
* No parameters

xbuf_51 
+ din1[51] din2[51] dout1[51] dout2[51] vdd vss 
+ dout_buf 
* No parameters

xbuf_52 
+ din1[52] din2[52] dout1[52] dout2[52] vdd vss 
+ dout_buf 
* No parameters

xbuf_53 
+ din1[53] din2[53] dout1[53] dout2[53] vdd vss 
+ dout_buf 
* No parameters

xbuf_54 
+ din1[54] din2[54] dout1[54] dout2[54] vdd vss 
+ dout_buf 
* No parameters

xbuf_55 
+ din1[55] din2[55] dout1[55] dout2[55] vdd vss 
+ dout_buf 
* No parameters

xbuf_56 
+ din1[56] din2[56] dout1[56] dout2[56] vdd vss 
+ dout_buf 
* No parameters

xbuf_57 
+ din1[57] din2[57] dout1[57] dout2[57] vdd vss 
+ dout_buf 
* No parameters

xbuf_58 
+ din1[58] din2[58] dout1[58] dout2[58] vdd vss 
+ dout_buf 
* No parameters

xbuf_59 
+ din1[59] din2[59] dout1[59] dout2[59] vdd vss 
+ dout_buf 
* No parameters

xbuf_60 
+ din1[60] din2[60] dout1[60] dout2[60] vdd vss 
+ dout_buf 
* No parameters

xbuf_61 
+ din1[61] din2[61] dout1[61] dout2[61] vdd vss 
+ dout_buf 
* No parameters

xbuf_62 
+ din1[62] din2[62] dout1[62] dout2[62] vdd vss 
+ dout_buf 
* No parameters

xbuf_63 
+ din1[63] din2[63] dout1[63] dout2[63] vdd vss 
+ dout_buf 
* No parameters

.ENDS

.SUBCKT we_control_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='8.0' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='12.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ we_control_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ we_control_and2_inv 
* No parameters

.ENDS

.SUBCKT we_control 
+ wr_en sel[1] sel[0] write_driver_en[1] write_driver_en[0] vdd vss 

xand2_0 
+ sel[0] wr_en write_driver_en[0] vdd vss 
+ we_control_and2 
* No parameters

xand2_1 
+ sel[1] wr_en write_driver_en[1] vdd vss 
+ we_control_and2 
* No parameters

.ENDS

.SUBCKT control_logic_delay_chain 
+ din dout vdd vss 

xinv_0 
+ din int[0] vdd vss 
+ control_logic_inv 
* No parameters

xinv_1 
+ int[0] int[1] vdd vss 
+ control_logic_inv 
* No parameters

xinv_2 
+ int[1] int[2] vdd vss 
+ control_logic_inv 
* No parameters

xinv_3 
+ int[2] int[3] vdd vss 
+ control_logic_inv 
* No parameters

xinv_4 
+ int[3] int[4] vdd vss 
+ control_logic_inv 
* No parameters

xinv_5 
+ int[4] int[5] vdd vss 
+ control_logic_inv 
* No parameters

xinv_6 
+ int[5] int[6] vdd vss 
+ control_logic_inv 
* No parameters

xinv_7 
+ int[6] int[7] vdd vss 
+ control_logic_inv 
* No parameters

xinv_8 
+ int[7] int[8] vdd vss 
+ control_logic_inv 
* No parameters

xinv_9 
+ int[8] int[9] vdd vss 
+ control_logic_inv 
* No parameters

xinv_10 
+ int[9] int[10] vdd vss 
+ control_logic_inv 
* No parameters

xinv_11 
+ int[10] int[11] vdd vss 
+ control_logic_inv 
* No parameters

xinv_12 
+ int[11] int[12] vdd vss 
+ control_logic_inv 
* No parameters

xinv_13 
+ int[12] int[13] vdd vss 
+ control_logic_inv 
* No parameters

xinv_14 
+ int[13] int[14] vdd vss 
+ control_logic_inv 
* No parameters

xinv_15 
+ int[14] int[15] vdd vss 
+ control_logic_inv 
* No parameters

xinv_16 
+ int[15] int[16] vdd vss 
+ control_logic_inv 
* No parameters

xinv_17 
+ int[16] int[17] vdd vss 
+ control_logic_inv 
* No parameters

xinv_18 
+ int[17] int[18] vdd vss 
+ control_logic_inv 
* No parameters

xinv_19 
+ int[18] int[19] vdd vss 
+ control_logic_inv 
* No parameters

xinv_20 
+ int[19] int[20] vdd vss 
+ control_logic_inv 
* No parameters

xinv_21 
+ int[20] int[21] vdd vss 
+ control_logic_inv 
* No parameters

xinv_22 
+ int[21] int[22] vdd vss 
+ control_logic_inv 
* No parameters

xinv_23 
+ int[22] int[23] vdd vss 
+ control_logic_inv 
* No parameters

xinv_24 
+ int[23] int[24] vdd vss 
+ control_logic_inv 
* No parameters

xinv_25 
+ int[24] int[25] vdd vss 
+ control_logic_inv 
* No parameters

xinv_26 
+ int[25] int[26] vdd vss 
+ control_logic_inv 
* No parameters

xinv_27 
+ int[26] int[27] vdd vss 
+ control_logic_inv 
* No parameters

xinv_28 
+ int[27] int[28] vdd vss 
+ control_logic_inv 
* No parameters

xinv_29 
+ int[28] int[29] vdd vss 
+ control_logic_inv 
* No parameters

xinv_30 
+ int[29] int[30] vdd vss 
+ control_logic_inv 
* No parameters

xinv_31 
+ int[30] int[31] vdd vss 
+ control_logic_inv 
* No parameters

xinv_32 
+ int[31] int[32] vdd vss 
+ control_logic_inv 
* No parameters

xinv_33 
+ int[32] int[33] vdd vss 
+ control_logic_inv 
* No parameters

xinv_34 
+ int[33] int[34] vdd vss 
+ control_logic_inv 
* No parameters

xinv_35 
+ int[34] int[35] vdd vss 
+ control_logic_inv 
* No parameters

xinv_36 
+ int[35] int[36] vdd vss 
+ control_logic_inv 
* No parameters

xinv_37 
+ int[36] int[37] vdd vss 
+ control_logic_inv 
* No parameters

xinv_38 
+ int[37] int[38] vdd vss 
+ control_logic_inv 
* No parameters

xinv_39 
+ int[38] int[39] vdd vss 
+ control_logic_inv 
* No parameters

xinv_40 
+ int[39] int[40] vdd vss 
+ control_logic_inv 
* No parameters

xinv_41 
+ int[40] int[41] vdd vss 
+ control_logic_inv 
* No parameters

xinv_42 
+ int[41] int[42] vdd vss 
+ control_logic_inv 
* No parameters

xinv_43 
+ int[42] int[43] vdd vss 
+ control_logic_inv 
* No parameters

xinv_44 
+ int[43] dout vdd vss 
+ control_logic_inv 
* No parameters

.ENDS

.SUBCKT sramgen_sram_128x64m2w64_replica_v1 
+ vdd vss clk din[63] din[62] din[61] din[60] din[59] din[58] din[57] din[56] din[55] din[54] din[53] din[52] din[51] din[50] din[49] din[48] din[47] din[46] din[45] din[44] din[43] din[42] din[41] din[40] din[39] din[38] din[37] din[36] din[35] din[34] din[33] din[32] din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] dout[63] dout[62] dout[61] dout[60] dout[59] dout[58] dout[57] dout[56] dout[55] dout[54] dout[53] dout[52] dout[51] dout[50] dout[49] dout[48] dout[47] dout[46] dout[45] dout[44] dout[43] dout[42] dout[41] dout[40] dout[39] dout[38] dout[37] dout[36] dout[35] dout[34] dout[33] dout[32] dout[31] dout[30] dout[29] dout[28] dout[27] dout[26] dout[25] dout[24] dout[23] dout[22] dout[21] dout[20] dout[19] dout[18] dout[17] dout[16] dout[15] dout[14] dout[13] dout[12] dout[11] dout[10] dout[9] dout[8] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] we addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] 

xdin_dffs 
+ vdd vss clk din[63] din[62] din[61] din[60] din[59] din[58] din[57] din[56] din[55] din[54] din[53] din[52] din[51] din[50] din[49] din[48] din[47] din[46] din[45] din[44] din[43] din[42] din[41] din[40] din[39] din[38] din[37] din[36] din[35] din[34] din[33] din[32] din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] bank_din[63] bank_din[62] bank_din[61] bank_din[60] bank_din[59] bank_din[58] bank_din[57] bank_din[56] bank_din[55] bank_din[54] bank_din[53] bank_din[52] bank_din[51] bank_din[50] bank_din[49] bank_din[48] bank_din[47] bank_din[46] bank_din[45] bank_din[44] bank_din[43] bank_din[42] bank_din[41] bank_din[40] bank_din[39] bank_din[38] bank_din[37] bank_din[36] bank_din[35] bank_din[34] bank_din[33] bank_din[32] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] dff_din_b[63] dff_din_b[62] dff_din_b[61] dff_din_b[60] dff_din_b[59] dff_din_b[58] dff_din_b[57] dff_din_b[56] dff_din_b[55] dff_din_b[54] dff_din_b[53] dff_din_b[52] dff_din_b[51] dff_din_b[50] dff_din_b[49] dff_din_b[48] dff_din_b[47] dff_din_b[46] dff_din_b[45] dff_din_b[44] dff_din_b[43] dff_din_b[42] dff_din_b[41] dff_din_b[40] dff_din_b[39] dff_din_b[38] dff_din_b[37] dff_din_b[36] dff_din_b[35] dff_din_b[34] dff_din_b[33] dff_din_b[32] dff_din_b[31] dff_din_b[30] dff_din_b[29] dff_din_b[28] dff_din_b[27] dff_din_b[26] dff_din_b[25] dff_din_b[24] dff_din_b[23] dff_din_b[22] dff_din_b[21] dff_din_b[20] dff_din_b[19] dff_din_b[18] dff_din_b[17] dff_din_b[16] dff_din_b[15] dff_din_b[14] dff_din_b[13] dff_din_b[12] dff_din_b[11] dff_din_b[10] dff_din_b[9] dff_din_b[8] dff_din_b[7] dff_din_b[6] dff_din_b[5] dff_din_b[4] dff_din_b[3] dff_din_b[2] dff_din_b[1] dff_din_b[0] 
+ data_dff_array 
* No parameters

xaddr_dffs 
+ vdd vss clk addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] bank_addr[6] bank_addr[5] bank_addr[4] bank_addr[3] bank_addr[2] bank_addr[1] bank_addr[0] bank_addr_b[6] bank_addr_b[5] bank_addr_b[4] bank_addr_b[3] bank_addr_b[2] bank_addr_b[1] bank_addr_b[0] 
+ addr_dff_array 
* No parameters

xwe_dff 
+ vdd vss clk we bank_we bank_we_b 
+ openram_dff 
* No parameters

xdecoder 
+ vdd vss bank_addr[6] bank_addr[5] bank_addr[4] bank_addr[3] bank_addr[2] bank_addr[1] bank_addr_b[6] bank_addr_b[5] bank_addr_b[4] bank_addr_b[3] bank_addr_b[2] bank_addr_b[1] wl_data[63] wl_data[62] wl_data[61] wl_data[60] wl_data[59] wl_data[58] wl_data[57] wl_data[56] wl_data[55] wl_data[54] wl_data[53] wl_data[52] wl_data[51] wl_data[50] wl_data[49] wl_data[48] wl_data[47] wl_data[46] wl_data[45] wl_data[44] wl_data[43] wl_data[42] wl_data[41] wl_data[40] wl_data[39] wl_data[38] wl_data[37] wl_data[36] wl_data[35] wl_data[34] wl_data[33] wl_data[32] wl_data[31] wl_data[30] wl_data[29] wl_data[28] wl_data[27] wl_data[26] wl_data[25] wl_data[24] wl_data[23] wl_data[22] wl_data[21] wl_data[20] wl_data[19] wl_data[18] wl_data[17] wl_data[16] wl_data[15] wl_data[14] wl_data[13] wl_data[12] wl_data[11] wl_data[10] wl_data[9] wl_data[8] wl_data[7] wl_data[6] wl_data[5] wl_data[4] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_data_b[63] wl_data_b[62] wl_data_b[61] wl_data_b[60] wl_data_b[59] wl_data_b[58] wl_data_b[57] wl_data_b[56] wl_data_b[55] wl_data_b[54] wl_data_b[53] wl_data_b[52] wl_data_b[51] wl_data_b[50] wl_data_b[49] wl_data_b[48] wl_data_b[47] wl_data_b[46] wl_data_b[45] wl_data_b[44] wl_data_b[43] wl_data_b[42] wl_data_b[41] wl_data_b[40] wl_data_b[39] wl_data_b[38] wl_data_b[37] wl_data_b[36] wl_data_b[35] wl_data_b[34] wl_data_b[33] wl_data_b[32] wl_data_b[31] wl_data_b[30] wl_data_b[29] wl_data_b[28] wl_data_b[27] wl_data_b[26] wl_data_b[25] wl_data_b[24] wl_data_b[23] wl_data_b[22] wl_data_b[21] wl_data_b[20] wl_data_b[19] wl_data_b[18] wl_data_b[17] wl_data_b[16] wl_data_b[15] wl_data_b[14] wl_data_b[13] wl_data_b[12] wl_data_b[11] wl_data_b[10] wl_data_b[9] wl_data_b[8] wl_data_b[7] wl_data_b[6] wl_data_b[5] wl_data_b[4] wl_data_b[3] wl_data_b[2] wl_data_b[1] wl_data_b[0] 
+ hierarchical_decoder 
* No parameters

xwl_driver_array 
+ vdd vss wl_data[63] wl_data[62] wl_data[61] wl_data[60] wl_data[59] wl_data[58] wl_data[57] wl_data[56] wl_data[55] wl_data[54] wl_data[53] wl_data[52] wl_data[51] wl_data[50] wl_data[49] wl_data[48] wl_data[47] wl_data[46] wl_data[45] wl_data[44] wl_data[43] wl_data[42] wl_data[41] wl_data[40] wl_data[39] wl_data[38] wl_data[37] wl_data[36] wl_data[35] wl_data[34] wl_data[33] wl_data[32] wl_data[31] wl_data[30] wl_data[29] wl_data[28] wl_data[27] wl_data[26] wl_data[25] wl_data[24] wl_data[23] wl_data[22] wl_data[21] wl_data[20] wl_data[19] wl_data[18] wl_data[17] wl_data[16] wl_data[15] wl_data[14] wl_data[13] wl_data[12] wl_data[11] wl_data[10] wl_data[9] wl_data[8] wl_data[7] wl_data[6] wl_data[5] wl_data[4] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_en wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] 
+ wordline_driver_array 
* No parameters

xbitcells 
+ vdd vss bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] vss vdd rbl rbr 
+ bitcell_array 
* No parameters

xprecharge_array 
+ vdd pc_b rbl bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0]  rbr br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0]  
+ precharge_array 
* No parameters

xwrite_mux_array 
+ write_driver_en[1] write_driver_en[0] bank_din[63] bank_din[62] bank_din[61] bank_din[60] bank_din[59] bank_din[58] bank_din[57] bank_din[56] bank_din[55] bank_din[54] bank_din[53] bank_din[52] bank_din[51] bank_din[50] bank_din[49] bank_din[48] bank_din[47] bank_din[46] bank_din[45] bank_din[44] bank_din[43] bank_din[42] bank_din[41] bank_din[40] bank_din[39] bank_din[38] bank_din[37] bank_din[36] bank_din[35] bank_din[34] bank_din[33] bank_din[32] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[63] bank_din_b[62] bank_din_b[61] bank_din_b[60] bank_din_b[59] bank_din_b[58] bank_din_b[57] bank_din_b[56] bank_din_b[55] bank_din_b[54] bank_din_b[53] bank_din_b[52] bank_din_b[51] bank_din_b[50] bank_din_b[49] bank_din_b[48] bank_din_b[47] bank_din_b[46] bank_din_b[45] bank_din_b[44] bank_din_b[43] bank_din_b[42] bank_din_b[41] bank_din_b[40] bank_din_b[39] bank_din_b[38] bank_din_b[37] bank_din_b[36] bank_din_b[35] bank_din_b[34] bank_din_b[33] bank_din_b[32] bank_din_b[31] bank_din_b[30] bank_din_b[29] bank_din_b[28] bank_din_b[27] bank_din_b[26] bank_din_b[25] bank_din_b[24] bank_din_b[23] bank_din_b[22] bank_din_b[21] bank_din_b[20] bank_din_b[19] bank_din_b[18] bank_din_b[17] bank_din_b[16] bank_din_b[15] bank_din_b[14] bank_din_b[13] bank_din_b[12] bank_din_b[11] bank_din_b[10] bank_din_b[9] bank_din_b[8] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 
+ write_mux_array 
* No parameters

xbank_addr_buf 
+ bank_addr[0] bank_addr_buf vdd vss 
+ control_logic_bufbuf_16 
* No parameters

xbank_addr_b_buf 
+ bank_addr_b[0] bank_addr_b_buf vdd vss 
+ control_logic_bufbuf_16 
* No parameters

xread_mux_array 
+ bank_addr_b_buf bank_addr_buf  bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_read[63] bl_read[62] bl_read[61] bl_read[60] bl_read[59] bl_read[58] bl_read[57] bl_read[56] bl_read[55] bl_read[54] bl_read[53] bl_read[52] bl_read[51] bl_read[50] bl_read[49] bl_read[48] bl_read[47] bl_read[46] bl_read[45] bl_read[44] bl_read[43] bl_read[42] bl_read[41] bl_read[40] bl_read[39] bl_read[38] bl_read[37] bl_read[36] bl_read[35] bl_read[34] bl_read[33] bl_read[32] bl_read[31] bl_read[30] bl_read[29] bl_read[28] bl_read[27] bl_read[26] bl_read[25] bl_read[24] bl_read[23] bl_read[22] bl_read[21] bl_read[20] bl_read[19] bl_read[18] bl_read[17] bl_read[16] bl_read[15] bl_read[14] bl_read[13] bl_read[12] bl_read[11] bl_read[10] bl_read[9] bl_read[8] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[63] br_read[62] br_read[61] br_read[60] br_read[59] br_read[58] br_read[57] br_read[56] br_read[55] br_read[54] br_read[53] br_read[52] br_read[51] br_read[50] br_read[49] br_read[48] br_read[47] br_read[46] br_read[45] br_read[44] br_read[43] br_read[42] br_read[41] br_read[40] br_read[39] br_read[38] br_read[37] br_read[36] br_read[35] br_read[34] br_read[33] br_read[32] br_read[31] br_read[30] br_read[29] br_read[28] br_read[27] br_read[26] br_read[25] br_read[24] br_read[23] br_read[22] br_read[21] br_read[20] br_read[19] br_read[18] br_read[17] br_read[16] br_read[15] br_read[14] br_read[13] br_read[12] br_read[11] br_read[10] br_read[9] br_read[8] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] vdd 
+ read_mux_array 
* No parameters

xcol_inv_array 
+ bank_din[63] bank_din[62] bank_din[61] bank_din[60] bank_din[59] bank_din[58] bank_din[57] bank_din[56] bank_din[55] bank_din[54] bank_din[53] bank_din[52] bank_din[51] bank_din[50] bank_din[49] bank_din[48] bank_din[47] bank_din[46] bank_din[45] bank_din[44] bank_din[43] bank_din[42] bank_din[41] bank_din[40] bank_din[39] bank_din[38] bank_din[37] bank_din[36] bank_din[35] bank_din[34] bank_din[33] bank_din[32] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[63] bank_din_b[62] bank_din_b[61] bank_din_b[60] bank_din_b[59] bank_din_b[58] bank_din_b[57] bank_din_b[56] bank_din_b[55] bank_din_b[54] bank_din_b[53] bank_din_b[52] bank_din_b[51] bank_din_b[50] bank_din_b[49] bank_din_b[48] bank_din_b[47] bank_din_b[46] bank_din_b[45] bank_din_b[44] bank_din_b[43] bank_din_b[42] bank_din_b[41] bank_din_b[40] bank_din_b[39] bank_din_b[38] bank_din_b[37] bank_din_b[36] bank_din_b[35] bank_din_b[34] bank_din_b[33] bank_din_b[32] bank_din_b[31] bank_din_b[30] bank_din_b[29] bank_din_b[28] bank_din_b[27] bank_din_b[26] bank_din_b[25] bank_din_b[24] bank_din_b[23] bank_din_b[22] bank_din_b[21] bank_din_b[20] bank_din_b[19] bank_din_b[18] bank_din_b[17] bank_din_b[16] bank_din_b[15] bank_din_b[14] bank_din_b[13] bank_din_b[12] bank_din_b[11] bank_din_b[10] bank_din_b[9] bank_din_b[8] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] vdd vss 
+ col_inv_array 
* No parameters

xsense_amp_array 
+ vdd vss sense_amp_en bl_read[63] bl_read[62] bl_read[61] bl_read[60] bl_read[59] bl_read[58] bl_read[57] bl_read[56] bl_read[55] bl_read[54] bl_read[53] bl_read[52] bl_read[51] bl_read[50] bl_read[49] bl_read[48] bl_read[47] bl_read[46] bl_read[45] bl_read[44] bl_read[43] bl_read[42] bl_read[41] bl_read[40] bl_read[39] bl_read[38] bl_read[37] bl_read[36] bl_read[35] bl_read[34] bl_read[33] bl_read[32] bl_read[31] bl_read[30] bl_read[29] bl_read[28] bl_read[27] bl_read[26] bl_read[25] bl_read[24] bl_read[23] bl_read[22] bl_read[21] bl_read[20] bl_read[19] bl_read[18] bl_read[17] bl_read[16] bl_read[15] bl_read[14] bl_read[13] bl_read[12] bl_read[11] bl_read[10] bl_read[9] bl_read[8] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[63] br_read[62] br_read[61] br_read[60] br_read[59] br_read[58] br_read[57] br_read[56] br_read[55] br_read[54] br_read[53] br_read[52] br_read[51] br_read[50] br_read[49] br_read[48] br_read[47] br_read[46] br_read[45] br_read[44] br_read[43] br_read[42] br_read[41] br_read[40] br_read[39] br_read[38] br_read[37] br_read[36] br_read[35] br_read[34] br_read[33] br_read[32] br_read[31] br_read[30] br_read[29] br_read[28] br_read[27] br_read[26] br_read[25] br_read[24] br_read[23] br_read[22] br_read[21] br_read[20] br_read[19] br_read[18] br_read[17] br_read[16] br_read[15] br_read[14] br_read[13] br_read[12] br_read[11] br_read[10] br_read[9] br_read[8] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] sa_outp[63] sa_outp[62] sa_outp[61] sa_outp[60] sa_outp[59] sa_outp[58] sa_outp[57] sa_outp[56] sa_outp[55] sa_outp[54] sa_outp[53] sa_outp[52] sa_outp[51] sa_outp[50] sa_outp[49] sa_outp[48] sa_outp[47] sa_outp[46] sa_outp[45] sa_outp[44] sa_outp[43] sa_outp[42] sa_outp[41] sa_outp[40] sa_outp[39] sa_outp[38] sa_outp[37] sa_outp[36] sa_outp[35] sa_outp[34] sa_outp[33] sa_outp[32] sa_outp[31] sa_outp[30] sa_outp[29] sa_outp[28] sa_outp[27] sa_outp[26] sa_outp[25] sa_outp[24] sa_outp[23] sa_outp[22] sa_outp[21] sa_outp[20] sa_outp[19] sa_outp[18] sa_outp[17] sa_outp[16] sa_outp[15] sa_outp[14] sa_outp[13] sa_outp[12] sa_outp[11] sa_outp[10] sa_outp[9] sa_outp[8] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[63] sa_outn[62] sa_outn[61] sa_outn[60] sa_outn[59] sa_outn[58] sa_outn[57] sa_outn[56] sa_outn[55] sa_outn[54] sa_outn[53] sa_outn[52] sa_outn[51] sa_outn[50] sa_outn[49] sa_outn[48] sa_outn[47] sa_outn[46] sa_outn[45] sa_outn[44] sa_outn[43] sa_outn[42] sa_outn[41] sa_outn[40] sa_outn[39] sa_outn[38] sa_outn[37] sa_outn[36] sa_outn[35] sa_outn[34] sa_outn[33] sa_outn[32] sa_outn[31] sa_outn[30] sa_outn[29] sa_outn[28] sa_outn[27] sa_outn[26] sa_outn[25] sa_outn[24] sa_outn[23] sa_outn[22] sa_outn[21] sa_outn[20] sa_outn[19] sa_outn[18] sa_outn[17] sa_outn[16] sa_outn[15] sa_outn[14] sa_outn[13] sa_outn[12] sa_outn[11] sa_outn[10] sa_outn[9] sa_outn[8] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] 
+ sense_amp_array 
* No parameters

xdout_buf_array 
+ sa_outp[63] sa_outp[62] sa_outp[61] sa_outp[60] sa_outp[59] sa_outp[58] sa_outp[57] sa_outp[56] sa_outp[55] sa_outp[54] sa_outp[53] sa_outp[52] sa_outp[51] sa_outp[50] sa_outp[49] sa_outp[48] sa_outp[47] sa_outp[46] sa_outp[45] sa_outp[44] sa_outp[43] sa_outp[42] sa_outp[41] sa_outp[40] sa_outp[39] sa_outp[38] sa_outp[37] sa_outp[36] sa_outp[35] sa_outp[34] sa_outp[33] sa_outp[32] sa_outp[31] sa_outp[30] sa_outp[29] sa_outp[28] sa_outp[27] sa_outp[26] sa_outp[25] sa_outp[24] sa_outp[23] sa_outp[22] sa_outp[21] sa_outp[20] sa_outp[19] sa_outp[18] sa_outp[17] sa_outp[16] sa_outp[15] sa_outp[14] sa_outp[13] sa_outp[12] sa_outp[11] sa_outp[10] sa_outp[9] sa_outp[8] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[63] sa_outn[62] sa_outn[61] sa_outn[60] sa_outn[59] sa_outn[58] sa_outn[57] sa_outn[56] sa_outn[55] sa_outn[54] sa_outn[53] sa_outn[52] sa_outn[51] sa_outn[50] sa_outn[49] sa_outn[48] sa_outn[47] sa_outn[46] sa_outn[45] sa_outn[44] sa_outn[43] sa_outn[42] sa_outn[41] sa_outn[40] sa_outn[39] sa_outn[38] sa_outn[37] sa_outn[36] sa_outn[35] sa_outn[34] sa_outn[33] sa_outn[32] sa_outn[31] sa_outn[30] sa_outn[29] sa_outn[28] sa_outn[27] sa_outn[26] sa_outn[25] sa_outn[24] sa_outn[23] sa_outn[22] sa_outn[21] sa_outn[20] sa_outn[19] sa_outn[18] sa_outn[17] sa_outn[16] sa_outn[15] sa_outn[14] sa_outn[13] sa_outn[12] sa_outn[11] sa_outn[10] sa_outn[9] sa_outn[8] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] dout[63] dout[62] dout[61] dout[60] dout[59] dout[58] dout[57] dout[56] dout[55] dout[54] dout[53] dout[52] dout[51] dout[50] dout[49] dout[48] dout[47] dout[46] dout[45] dout[44] dout[43] dout[42] dout[41] dout[40] dout[39] dout[38] dout[37] dout[36] dout[35] dout[34] dout[33] dout[32] dout[31] dout[30] dout[29] dout[28] dout[27] dout[26] dout[25] dout[24] dout[23] dout[22] dout[21] dout[20] dout[19] dout[18] dout[17] dout[16] dout[15] dout[14] dout[13] dout[12] dout[11] dout[10] dout[9] dout[8] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] dout_b[63] dout_b[62] dout_b[61] dout_b[60] dout_b[59] dout_b[58] dout_b[57] dout_b[56] dout_b[55] dout_b[54] dout_b[53] dout_b[52] dout_b[51] dout_b[50] dout_b[49] dout_b[48] dout_b[47] dout_b[46] dout_b[45] dout_b[44] dout_b[43] dout_b[42] dout_b[41] dout_b[40] dout_b[39] dout_b[38] dout_b[37] dout_b[36] dout_b[35] dout_b[34] dout_b[33] dout_b[32] dout_b[31] dout_b[30] dout_b[29] dout_b[28] dout_b[27] dout_b[26] dout_b[25] dout_b[24] dout_b[23] dout_b[22] dout_b[21] dout_b[20] dout_b[19] dout_b[18] dout_b[17] dout_b[16] dout_b[15] dout_b[14] dout_b[13] dout_b[12] dout_b[11] dout_b[10] dout_b[9] dout_b[8] dout_b[7] dout_b[6] dout_b[5] dout_b[4] dout_b[3] dout_b[2] dout_b[1] dout_b[0] vdd vss 
+ dout_buf_array 
* No parameters

xcontrol_logic 
+ clk bank_we rbl pc_b wl_en wr_en sense_amp_en vdd vss 
+ sramgen_control_replica_v1 
* No parameters

xwe_control 
+ wr_en bank_addr[0] bank_addr_b[0]  write_driver_en[1] write_driver_en[0] vdd vss 
+ we_control 
* No parameters

.ENDS

